`include "Decoder_Parameters.v"
module get_msgini(
    input clk,
    input rst_n,
    input [`Zc*`VWidth-1:0] data_in, //输入目的是分割一个方阵的元素为Zc/DPU_num组
    input [`APP_addr_width-2:0] addr_in,
	input en_in,
    output reg [`inNum*`VWidth-1:0] data_out //输出32长度，就是DPU并行度的长度
	// output reg [`APP_addr_width-2:0] addr_out
);

reg [`APP_addr_width-2:0] addr_in_D0;
// always @(posedge clk or negedge rst_n)
// begin
// 	if(!rst_n)
// 	begin
// 		addr_out <= 0;
// 	end
// 	else
// 	begin
// 		addr_out <= addr_in;
// 	end
// end

always @(posedge clk or negedge rst_n)
begin
	if(!rst_n)
	begin
		addr_in_D0 <= 0;
	end
	else
	begin
		addr_in_D0 <= addr_in;
	end
end

always @(posedge clk or negedge rst_n)
begin
	if(!rst_n)
	begin
		data_out <= 0;
	end
	else if(en_in)
	begin
		case(addr_in)
			0:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+1)-1:`VWidth*(`APPRam_depth*31+0)],data_in[`VWidth*(`APPRam_depth*30+1)-1:`VWidth*(`APPRam_depth*30+0)],data_in[`VWidth*(`APPRam_depth*29+1)-1:`VWidth*(`APPRam_depth*29+0)],data_in[`VWidth*(`APPRam_depth*28+1)-1:`VWidth*(`APPRam_depth*28+0)],data_in[`VWidth*(`APPRam_depth*27+1)-1:`VWidth*(`APPRam_depth*27+0)],data_in[`VWidth*(`APPRam_depth*26+1)-1:`VWidth*(`APPRam_depth*26+0)],data_in[`VWidth*(`APPRam_depth*25+1)-1:`VWidth*(`APPRam_depth*25+0)],data_in[`VWidth*(`APPRam_depth*24+1)-1:`VWidth*(`APPRam_depth*24+0)],data_in[`VWidth*(`APPRam_depth*23+1)-1:`VWidth*(`APPRam_depth*23+0)],data_in[`VWidth*(`APPRam_depth*22+1)-1:`VWidth*(`APPRam_depth*22+0)],data_in[`VWidth*(`APPRam_depth*21+1)-1:`VWidth*(`APPRam_depth*21+0)],data_in[`VWidth*(`APPRam_depth*20+1)-1:`VWidth*(`APPRam_depth*20+0)],data_in[`VWidth*(`APPRam_depth*19+1)-1:`VWidth*(`APPRam_depth*19+0)],data_in[`VWidth*(`APPRam_depth*18+1)-1:`VWidth*(`APPRam_depth*18+0)],data_in[`VWidth*(`APPRam_depth*17+1)-1:`VWidth*(`APPRam_depth*17+0)],data_in[`VWidth*(`APPRam_depth*16+1)-1:`VWidth*(`APPRam_depth*16+0)],data_in[`VWidth*(`APPRam_depth*15+1)-1:`VWidth*(`APPRam_depth*15+0)],data_in[`VWidth*(`APPRam_depth*14+1)-1:`VWidth*(`APPRam_depth*14+0)],data_in[`VWidth*(`APPRam_depth*13+1)-1:`VWidth*(`APPRam_depth*13+0)],data_in[`VWidth*(`APPRam_depth*12+1)-1:`VWidth*(`APPRam_depth*12+0)],data_in[`VWidth*(`APPRam_depth*11+1)-1:`VWidth*(`APPRam_depth*11+0)],data_in[`VWidth*(`APPRam_depth*10+1)-1:`VWidth*(`APPRam_depth*10+0)],data_in[`VWidth*(`APPRam_depth*9+1)-1:`VWidth*(`APPRam_depth*9+0)],data_in[`VWidth*(`APPRam_depth*8+1)-1:`VWidth*(`APPRam_depth*8+0)],data_in[`VWidth*(`APPRam_depth*7+1)-1:`VWidth*(`APPRam_depth*7+0)],data_in[`VWidth*(`APPRam_depth*6+1)-1:`VWidth*(`APPRam_depth*6+0)],data_in[`VWidth*(`APPRam_depth*5+1)-1:`VWidth*(`APPRam_depth*5+0)],data_in[`VWidth*(`APPRam_depth*4+1)-1:`VWidth*(`APPRam_depth*4+0)],data_in[`VWidth*(`APPRam_depth*3+1)-1:`VWidth*(`APPRam_depth*3+0)],data_in[`VWidth*(`APPRam_depth*2+1)-1:`VWidth*(`APPRam_depth*2+0)],data_in[`VWidth*(`APPRam_depth*1+1)-1:`VWidth*(`APPRam_depth*1+0)],data_in[`VWidth*(`APPRam_depth*0+1)-1:`VWidth*(`APPRam_depth*0+0)]};
			end
			1:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+2)-1:`VWidth*(`APPRam_depth*31+1)],data_in[`VWidth*(`APPRam_depth*30+2)-1:`VWidth*(`APPRam_depth*30+1)],data_in[`VWidth*(`APPRam_depth*29+2)-1:`VWidth*(`APPRam_depth*29+1)],data_in[`VWidth*(`APPRam_depth*28+2)-1:`VWidth*(`APPRam_depth*28+1)],data_in[`VWidth*(`APPRam_depth*27+2)-1:`VWidth*(`APPRam_depth*27+1)],data_in[`VWidth*(`APPRam_depth*26+2)-1:`VWidth*(`APPRam_depth*26+1)],data_in[`VWidth*(`APPRam_depth*25+2)-1:`VWidth*(`APPRam_depth*25+1)],data_in[`VWidth*(`APPRam_depth*24+2)-1:`VWidth*(`APPRam_depth*24+1)],data_in[`VWidth*(`APPRam_depth*23+2)-1:`VWidth*(`APPRam_depth*23+1)],data_in[`VWidth*(`APPRam_depth*22+2)-1:`VWidth*(`APPRam_depth*22+1)],data_in[`VWidth*(`APPRam_depth*21+2)-1:`VWidth*(`APPRam_depth*21+1)],data_in[`VWidth*(`APPRam_depth*20+2)-1:`VWidth*(`APPRam_depth*20+1)],data_in[`VWidth*(`APPRam_depth*19+2)-1:`VWidth*(`APPRam_depth*19+1)],data_in[`VWidth*(`APPRam_depth*18+2)-1:`VWidth*(`APPRam_depth*18+1)],data_in[`VWidth*(`APPRam_depth*17+2)-1:`VWidth*(`APPRam_depth*17+1)],data_in[`VWidth*(`APPRam_depth*16+2)-1:`VWidth*(`APPRam_depth*16+1)],data_in[`VWidth*(`APPRam_depth*15+2)-1:`VWidth*(`APPRam_depth*15+1)],data_in[`VWidth*(`APPRam_depth*14+2)-1:`VWidth*(`APPRam_depth*14+1)],data_in[`VWidth*(`APPRam_depth*13+2)-1:`VWidth*(`APPRam_depth*13+1)],data_in[`VWidth*(`APPRam_depth*12+2)-1:`VWidth*(`APPRam_depth*12+1)],data_in[`VWidth*(`APPRam_depth*11+2)-1:`VWidth*(`APPRam_depth*11+1)],data_in[`VWidth*(`APPRam_depth*10+2)-1:`VWidth*(`APPRam_depth*10+1)],data_in[`VWidth*(`APPRam_depth*9+2)-1:`VWidth*(`APPRam_depth*9+1)],data_in[`VWidth*(`APPRam_depth*8+2)-1:`VWidth*(`APPRam_depth*8+1)],data_in[`VWidth*(`APPRam_depth*7+2)-1:`VWidth*(`APPRam_depth*7+1)],data_in[`VWidth*(`APPRam_depth*6+2)-1:`VWidth*(`APPRam_depth*6+1)],data_in[`VWidth*(`APPRam_depth*5+2)-1:`VWidth*(`APPRam_depth*5+1)],data_in[`VWidth*(`APPRam_depth*4+2)-1:`VWidth*(`APPRam_depth*4+1)],data_in[`VWidth*(`APPRam_depth*3+2)-1:`VWidth*(`APPRam_depth*3+1)],data_in[`VWidth*(`APPRam_depth*2+2)-1:`VWidth*(`APPRam_depth*2+1)],data_in[`VWidth*(`APPRam_depth*1+2)-1:`VWidth*(`APPRam_depth*1+1)],data_in[`VWidth*(`APPRam_depth*0+2)-1:`VWidth*(`APPRam_depth*0+1)]};
			end
			2:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+3)-1:`VWidth*(`APPRam_depth*31+2)],data_in[`VWidth*(`APPRam_depth*30+3)-1:`VWidth*(`APPRam_depth*30+2)],data_in[`VWidth*(`APPRam_depth*29+3)-1:`VWidth*(`APPRam_depth*29+2)],data_in[`VWidth*(`APPRam_depth*28+3)-1:`VWidth*(`APPRam_depth*28+2)],data_in[`VWidth*(`APPRam_depth*27+3)-1:`VWidth*(`APPRam_depth*27+2)],data_in[`VWidth*(`APPRam_depth*26+3)-1:`VWidth*(`APPRam_depth*26+2)],data_in[`VWidth*(`APPRam_depth*25+3)-1:`VWidth*(`APPRam_depth*25+2)],data_in[`VWidth*(`APPRam_depth*24+3)-1:`VWidth*(`APPRam_depth*24+2)],data_in[`VWidth*(`APPRam_depth*23+3)-1:`VWidth*(`APPRam_depth*23+2)],data_in[`VWidth*(`APPRam_depth*22+3)-1:`VWidth*(`APPRam_depth*22+2)],data_in[`VWidth*(`APPRam_depth*21+3)-1:`VWidth*(`APPRam_depth*21+2)],data_in[`VWidth*(`APPRam_depth*20+3)-1:`VWidth*(`APPRam_depth*20+2)],data_in[`VWidth*(`APPRam_depth*19+3)-1:`VWidth*(`APPRam_depth*19+2)],data_in[`VWidth*(`APPRam_depth*18+3)-1:`VWidth*(`APPRam_depth*18+2)],data_in[`VWidth*(`APPRam_depth*17+3)-1:`VWidth*(`APPRam_depth*17+2)],data_in[`VWidth*(`APPRam_depth*16+3)-1:`VWidth*(`APPRam_depth*16+2)],data_in[`VWidth*(`APPRam_depth*15+3)-1:`VWidth*(`APPRam_depth*15+2)],data_in[`VWidth*(`APPRam_depth*14+3)-1:`VWidth*(`APPRam_depth*14+2)],data_in[`VWidth*(`APPRam_depth*13+3)-1:`VWidth*(`APPRam_depth*13+2)],data_in[`VWidth*(`APPRam_depth*12+3)-1:`VWidth*(`APPRam_depth*12+2)],data_in[`VWidth*(`APPRam_depth*11+3)-1:`VWidth*(`APPRam_depth*11+2)],data_in[`VWidth*(`APPRam_depth*10+3)-1:`VWidth*(`APPRam_depth*10+2)],data_in[`VWidth*(`APPRam_depth*9+3)-1:`VWidth*(`APPRam_depth*9+2)],data_in[`VWidth*(`APPRam_depth*8+3)-1:`VWidth*(`APPRam_depth*8+2)],data_in[`VWidth*(`APPRam_depth*7+3)-1:`VWidth*(`APPRam_depth*7+2)],data_in[`VWidth*(`APPRam_depth*6+3)-1:`VWidth*(`APPRam_depth*6+2)],data_in[`VWidth*(`APPRam_depth*5+3)-1:`VWidth*(`APPRam_depth*5+2)],data_in[`VWidth*(`APPRam_depth*4+3)-1:`VWidth*(`APPRam_depth*4+2)],data_in[`VWidth*(`APPRam_depth*3+3)-1:`VWidth*(`APPRam_depth*3+2)],data_in[`VWidth*(`APPRam_depth*2+3)-1:`VWidth*(`APPRam_depth*2+2)],data_in[`VWidth*(`APPRam_depth*1+3)-1:`VWidth*(`APPRam_depth*1+2)],data_in[`VWidth*(`APPRam_depth*0+3)-1:`VWidth*(`APPRam_depth*0+2)]};
			end
			3:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+4)-1:`VWidth*(`APPRam_depth*31+3)],data_in[`VWidth*(`APPRam_depth*30+4)-1:`VWidth*(`APPRam_depth*30+3)],data_in[`VWidth*(`APPRam_depth*29+4)-1:`VWidth*(`APPRam_depth*29+3)],data_in[`VWidth*(`APPRam_depth*28+4)-1:`VWidth*(`APPRam_depth*28+3)],data_in[`VWidth*(`APPRam_depth*27+4)-1:`VWidth*(`APPRam_depth*27+3)],data_in[`VWidth*(`APPRam_depth*26+4)-1:`VWidth*(`APPRam_depth*26+3)],data_in[`VWidth*(`APPRam_depth*25+4)-1:`VWidth*(`APPRam_depth*25+3)],data_in[`VWidth*(`APPRam_depth*24+4)-1:`VWidth*(`APPRam_depth*24+3)],data_in[`VWidth*(`APPRam_depth*23+4)-1:`VWidth*(`APPRam_depth*23+3)],data_in[`VWidth*(`APPRam_depth*22+4)-1:`VWidth*(`APPRam_depth*22+3)],data_in[`VWidth*(`APPRam_depth*21+4)-1:`VWidth*(`APPRam_depth*21+3)],data_in[`VWidth*(`APPRam_depth*20+4)-1:`VWidth*(`APPRam_depth*20+3)],data_in[`VWidth*(`APPRam_depth*19+4)-1:`VWidth*(`APPRam_depth*19+3)],data_in[`VWidth*(`APPRam_depth*18+4)-1:`VWidth*(`APPRam_depth*18+3)],data_in[`VWidth*(`APPRam_depth*17+4)-1:`VWidth*(`APPRam_depth*17+3)],data_in[`VWidth*(`APPRam_depth*16+4)-1:`VWidth*(`APPRam_depth*16+3)],data_in[`VWidth*(`APPRam_depth*15+4)-1:`VWidth*(`APPRam_depth*15+3)],data_in[`VWidth*(`APPRam_depth*14+4)-1:`VWidth*(`APPRam_depth*14+3)],data_in[`VWidth*(`APPRam_depth*13+4)-1:`VWidth*(`APPRam_depth*13+3)],data_in[`VWidth*(`APPRam_depth*12+4)-1:`VWidth*(`APPRam_depth*12+3)],data_in[`VWidth*(`APPRam_depth*11+4)-1:`VWidth*(`APPRam_depth*11+3)],data_in[`VWidth*(`APPRam_depth*10+4)-1:`VWidth*(`APPRam_depth*10+3)],data_in[`VWidth*(`APPRam_depth*9+4)-1:`VWidth*(`APPRam_depth*9+3)],data_in[`VWidth*(`APPRam_depth*8+4)-1:`VWidth*(`APPRam_depth*8+3)],data_in[`VWidth*(`APPRam_depth*7+4)-1:`VWidth*(`APPRam_depth*7+3)],data_in[`VWidth*(`APPRam_depth*6+4)-1:`VWidth*(`APPRam_depth*6+3)],data_in[`VWidth*(`APPRam_depth*5+4)-1:`VWidth*(`APPRam_depth*5+3)],data_in[`VWidth*(`APPRam_depth*4+4)-1:`VWidth*(`APPRam_depth*4+3)],data_in[`VWidth*(`APPRam_depth*3+4)-1:`VWidth*(`APPRam_depth*3+3)],data_in[`VWidth*(`APPRam_depth*2+4)-1:`VWidth*(`APPRam_depth*2+3)],data_in[`VWidth*(`APPRam_depth*1+4)-1:`VWidth*(`APPRam_depth*1+3)],data_in[`VWidth*(`APPRam_depth*0+4)-1:`VWidth*(`APPRam_depth*0+3)]};
			end
			4:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+5)-1:`VWidth*(`APPRam_depth*31+4)],data_in[`VWidth*(`APPRam_depth*30+5)-1:`VWidth*(`APPRam_depth*30+4)],data_in[`VWidth*(`APPRam_depth*29+5)-1:`VWidth*(`APPRam_depth*29+4)],data_in[`VWidth*(`APPRam_depth*28+5)-1:`VWidth*(`APPRam_depth*28+4)],data_in[`VWidth*(`APPRam_depth*27+5)-1:`VWidth*(`APPRam_depth*27+4)],data_in[`VWidth*(`APPRam_depth*26+5)-1:`VWidth*(`APPRam_depth*26+4)],data_in[`VWidth*(`APPRam_depth*25+5)-1:`VWidth*(`APPRam_depth*25+4)],data_in[`VWidth*(`APPRam_depth*24+5)-1:`VWidth*(`APPRam_depth*24+4)],data_in[`VWidth*(`APPRam_depth*23+5)-1:`VWidth*(`APPRam_depth*23+4)],data_in[`VWidth*(`APPRam_depth*22+5)-1:`VWidth*(`APPRam_depth*22+4)],data_in[`VWidth*(`APPRam_depth*21+5)-1:`VWidth*(`APPRam_depth*21+4)],data_in[`VWidth*(`APPRam_depth*20+5)-1:`VWidth*(`APPRam_depth*20+4)],data_in[`VWidth*(`APPRam_depth*19+5)-1:`VWidth*(`APPRam_depth*19+4)],data_in[`VWidth*(`APPRam_depth*18+5)-1:`VWidth*(`APPRam_depth*18+4)],data_in[`VWidth*(`APPRam_depth*17+5)-1:`VWidth*(`APPRam_depth*17+4)],data_in[`VWidth*(`APPRam_depth*16+5)-1:`VWidth*(`APPRam_depth*16+4)],data_in[`VWidth*(`APPRam_depth*15+5)-1:`VWidth*(`APPRam_depth*15+4)],data_in[`VWidth*(`APPRam_depth*14+5)-1:`VWidth*(`APPRam_depth*14+4)],data_in[`VWidth*(`APPRam_depth*13+5)-1:`VWidth*(`APPRam_depth*13+4)],data_in[`VWidth*(`APPRam_depth*12+5)-1:`VWidth*(`APPRam_depth*12+4)],data_in[`VWidth*(`APPRam_depth*11+5)-1:`VWidth*(`APPRam_depth*11+4)],data_in[`VWidth*(`APPRam_depth*10+5)-1:`VWidth*(`APPRam_depth*10+4)],data_in[`VWidth*(`APPRam_depth*9+5)-1:`VWidth*(`APPRam_depth*9+4)],data_in[`VWidth*(`APPRam_depth*8+5)-1:`VWidth*(`APPRam_depth*8+4)],data_in[`VWidth*(`APPRam_depth*7+5)-1:`VWidth*(`APPRam_depth*7+4)],data_in[`VWidth*(`APPRam_depth*6+5)-1:`VWidth*(`APPRam_depth*6+4)],data_in[`VWidth*(`APPRam_depth*5+5)-1:`VWidth*(`APPRam_depth*5+4)],data_in[`VWidth*(`APPRam_depth*4+5)-1:`VWidth*(`APPRam_depth*4+4)],data_in[`VWidth*(`APPRam_depth*3+5)-1:`VWidth*(`APPRam_depth*3+4)],data_in[`VWidth*(`APPRam_depth*2+5)-1:`VWidth*(`APPRam_depth*2+4)],data_in[`VWidth*(`APPRam_depth*1+5)-1:`VWidth*(`APPRam_depth*1+4)],data_in[`VWidth*(`APPRam_depth*0+5)-1:`VWidth*(`APPRam_depth*0+4)]};
			end
			5:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+6)-1:`VWidth*(`APPRam_depth*31+5)],data_in[`VWidth*(`APPRam_depth*30+6)-1:`VWidth*(`APPRam_depth*30+5)],data_in[`VWidth*(`APPRam_depth*29+6)-1:`VWidth*(`APPRam_depth*29+5)],data_in[`VWidth*(`APPRam_depth*28+6)-1:`VWidth*(`APPRam_depth*28+5)],data_in[`VWidth*(`APPRam_depth*27+6)-1:`VWidth*(`APPRam_depth*27+5)],data_in[`VWidth*(`APPRam_depth*26+6)-1:`VWidth*(`APPRam_depth*26+5)],data_in[`VWidth*(`APPRam_depth*25+6)-1:`VWidth*(`APPRam_depth*25+5)],data_in[`VWidth*(`APPRam_depth*24+6)-1:`VWidth*(`APPRam_depth*24+5)],data_in[`VWidth*(`APPRam_depth*23+6)-1:`VWidth*(`APPRam_depth*23+5)],data_in[`VWidth*(`APPRam_depth*22+6)-1:`VWidth*(`APPRam_depth*22+5)],data_in[`VWidth*(`APPRam_depth*21+6)-1:`VWidth*(`APPRam_depth*21+5)],data_in[`VWidth*(`APPRam_depth*20+6)-1:`VWidth*(`APPRam_depth*20+5)],data_in[`VWidth*(`APPRam_depth*19+6)-1:`VWidth*(`APPRam_depth*19+5)],data_in[`VWidth*(`APPRam_depth*18+6)-1:`VWidth*(`APPRam_depth*18+5)],data_in[`VWidth*(`APPRam_depth*17+6)-1:`VWidth*(`APPRam_depth*17+5)],data_in[`VWidth*(`APPRam_depth*16+6)-1:`VWidth*(`APPRam_depth*16+5)],data_in[`VWidth*(`APPRam_depth*15+6)-1:`VWidth*(`APPRam_depth*15+5)],data_in[`VWidth*(`APPRam_depth*14+6)-1:`VWidth*(`APPRam_depth*14+5)],data_in[`VWidth*(`APPRam_depth*13+6)-1:`VWidth*(`APPRam_depth*13+5)],data_in[`VWidth*(`APPRam_depth*12+6)-1:`VWidth*(`APPRam_depth*12+5)],data_in[`VWidth*(`APPRam_depth*11+6)-1:`VWidth*(`APPRam_depth*11+5)],data_in[`VWidth*(`APPRam_depth*10+6)-1:`VWidth*(`APPRam_depth*10+5)],data_in[`VWidth*(`APPRam_depth*9+6)-1:`VWidth*(`APPRam_depth*9+5)],data_in[`VWidth*(`APPRam_depth*8+6)-1:`VWidth*(`APPRam_depth*8+5)],data_in[`VWidth*(`APPRam_depth*7+6)-1:`VWidth*(`APPRam_depth*7+5)],data_in[`VWidth*(`APPRam_depth*6+6)-1:`VWidth*(`APPRam_depth*6+5)],data_in[`VWidth*(`APPRam_depth*5+6)-1:`VWidth*(`APPRam_depth*5+5)],data_in[`VWidth*(`APPRam_depth*4+6)-1:`VWidth*(`APPRam_depth*4+5)],data_in[`VWidth*(`APPRam_depth*3+6)-1:`VWidth*(`APPRam_depth*3+5)],data_in[`VWidth*(`APPRam_depth*2+6)-1:`VWidth*(`APPRam_depth*2+5)],data_in[`VWidth*(`APPRam_depth*1+6)-1:`VWidth*(`APPRam_depth*1+5)],data_in[`VWidth*(`APPRam_depth*0+6)-1:`VWidth*(`APPRam_depth*0+5)]};
			end
			6:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+7)-1:`VWidth*(`APPRam_depth*31+6)],data_in[`VWidth*(`APPRam_depth*30+7)-1:`VWidth*(`APPRam_depth*30+6)],data_in[`VWidth*(`APPRam_depth*29+7)-1:`VWidth*(`APPRam_depth*29+6)],data_in[`VWidth*(`APPRam_depth*28+7)-1:`VWidth*(`APPRam_depth*28+6)],data_in[`VWidth*(`APPRam_depth*27+7)-1:`VWidth*(`APPRam_depth*27+6)],data_in[`VWidth*(`APPRam_depth*26+7)-1:`VWidth*(`APPRam_depth*26+6)],data_in[`VWidth*(`APPRam_depth*25+7)-1:`VWidth*(`APPRam_depth*25+6)],data_in[`VWidth*(`APPRam_depth*24+7)-1:`VWidth*(`APPRam_depth*24+6)],data_in[`VWidth*(`APPRam_depth*23+7)-1:`VWidth*(`APPRam_depth*23+6)],data_in[`VWidth*(`APPRam_depth*22+7)-1:`VWidth*(`APPRam_depth*22+6)],data_in[`VWidth*(`APPRam_depth*21+7)-1:`VWidth*(`APPRam_depth*21+6)],data_in[`VWidth*(`APPRam_depth*20+7)-1:`VWidth*(`APPRam_depth*20+6)],data_in[`VWidth*(`APPRam_depth*19+7)-1:`VWidth*(`APPRam_depth*19+6)],data_in[`VWidth*(`APPRam_depth*18+7)-1:`VWidth*(`APPRam_depth*18+6)],data_in[`VWidth*(`APPRam_depth*17+7)-1:`VWidth*(`APPRam_depth*17+6)],data_in[`VWidth*(`APPRam_depth*16+7)-1:`VWidth*(`APPRam_depth*16+6)],data_in[`VWidth*(`APPRam_depth*15+7)-1:`VWidth*(`APPRam_depth*15+6)],data_in[`VWidth*(`APPRam_depth*14+7)-1:`VWidth*(`APPRam_depth*14+6)],data_in[`VWidth*(`APPRam_depth*13+7)-1:`VWidth*(`APPRam_depth*13+6)],data_in[`VWidth*(`APPRam_depth*12+7)-1:`VWidth*(`APPRam_depth*12+6)],data_in[`VWidth*(`APPRam_depth*11+7)-1:`VWidth*(`APPRam_depth*11+6)],data_in[`VWidth*(`APPRam_depth*10+7)-1:`VWidth*(`APPRam_depth*10+6)],data_in[`VWidth*(`APPRam_depth*9+7)-1:`VWidth*(`APPRam_depth*9+6)],data_in[`VWidth*(`APPRam_depth*8+7)-1:`VWidth*(`APPRam_depth*8+6)],data_in[`VWidth*(`APPRam_depth*7+7)-1:`VWidth*(`APPRam_depth*7+6)],data_in[`VWidth*(`APPRam_depth*6+7)-1:`VWidth*(`APPRam_depth*6+6)],data_in[`VWidth*(`APPRam_depth*5+7)-1:`VWidth*(`APPRam_depth*5+6)],data_in[`VWidth*(`APPRam_depth*4+7)-1:`VWidth*(`APPRam_depth*4+6)],data_in[`VWidth*(`APPRam_depth*3+7)-1:`VWidth*(`APPRam_depth*3+6)],data_in[`VWidth*(`APPRam_depth*2+7)-1:`VWidth*(`APPRam_depth*2+6)],data_in[`VWidth*(`APPRam_depth*1+7)-1:`VWidth*(`APPRam_depth*1+6)],data_in[`VWidth*(`APPRam_depth*0+7)-1:`VWidth*(`APPRam_depth*0+6)]};
			end
			7:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+8)-1:`VWidth*(`APPRam_depth*31+7)],data_in[`VWidth*(`APPRam_depth*30+8)-1:`VWidth*(`APPRam_depth*30+7)],data_in[`VWidth*(`APPRam_depth*29+8)-1:`VWidth*(`APPRam_depth*29+7)],data_in[`VWidth*(`APPRam_depth*28+8)-1:`VWidth*(`APPRam_depth*28+7)],data_in[`VWidth*(`APPRam_depth*27+8)-1:`VWidth*(`APPRam_depth*27+7)],data_in[`VWidth*(`APPRam_depth*26+8)-1:`VWidth*(`APPRam_depth*26+7)],data_in[`VWidth*(`APPRam_depth*25+8)-1:`VWidth*(`APPRam_depth*25+7)],data_in[`VWidth*(`APPRam_depth*24+8)-1:`VWidth*(`APPRam_depth*24+7)],data_in[`VWidth*(`APPRam_depth*23+8)-1:`VWidth*(`APPRam_depth*23+7)],data_in[`VWidth*(`APPRam_depth*22+8)-1:`VWidth*(`APPRam_depth*22+7)],data_in[`VWidth*(`APPRam_depth*21+8)-1:`VWidth*(`APPRam_depth*21+7)],data_in[`VWidth*(`APPRam_depth*20+8)-1:`VWidth*(`APPRam_depth*20+7)],data_in[`VWidth*(`APPRam_depth*19+8)-1:`VWidth*(`APPRam_depth*19+7)],data_in[`VWidth*(`APPRam_depth*18+8)-1:`VWidth*(`APPRam_depth*18+7)],data_in[`VWidth*(`APPRam_depth*17+8)-1:`VWidth*(`APPRam_depth*17+7)],data_in[`VWidth*(`APPRam_depth*16+8)-1:`VWidth*(`APPRam_depth*16+7)],data_in[`VWidth*(`APPRam_depth*15+8)-1:`VWidth*(`APPRam_depth*15+7)],data_in[`VWidth*(`APPRam_depth*14+8)-1:`VWidth*(`APPRam_depth*14+7)],data_in[`VWidth*(`APPRam_depth*13+8)-1:`VWidth*(`APPRam_depth*13+7)],data_in[`VWidth*(`APPRam_depth*12+8)-1:`VWidth*(`APPRam_depth*12+7)],data_in[`VWidth*(`APPRam_depth*11+8)-1:`VWidth*(`APPRam_depth*11+7)],data_in[`VWidth*(`APPRam_depth*10+8)-1:`VWidth*(`APPRam_depth*10+7)],data_in[`VWidth*(`APPRam_depth*9+8)-1:`VWidth*(`APPRam_depth*9+7)],data_in[`VWidth*(`APPRam_depth*8+8)-1:`VWidth*(`APPRam_depth*8+7)],data_in[`VWidth*(`APPRam_depth*7+8)-1:`VWidth*(`APPRam_depth*7+7)],data_in[`VWidth*(`APPRam_depth*6+8)-1:`VWidth*(`APPRam_depth*6+7)],data_in[`VWidth*(`APPRam_depth*5+8)-1:`VWidth*(`APPRam_depth*5+7)],data_in[`VWidth*(`APPRam_depth*4+8)-1:`VWidth*(`APPRam_depth*4+7)],data_in[`VWidth*(`APPRam_depth*3+8)-1:`VWidth*(`APPRam_depth*3+7)],data_in[`VWidth*(`APPRam_depth*2+8)-1:`VWidth*(`APPRam_depth*2+7)],data_in[`VWidth*(`APPRam_depth*1+8)-1:`VWidth*(`APPRam_depth*1+7)],data_in[`VWidth*(`APPRam_depth*0+8)-1:`VWidth*(`APPRam_depth*0+7)]};
			end
			8:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+9)-1:`VWidth*(`APPRam_depth*31+8)],data_in[`VWidth*(`APPRam_depth*30+9)-1:`VWidth*(`APPRam_depth*30+8)],data_in[`VWidth*(`APPRam_depth*29+9)-1:`VWidth*(`APPRam_depth*29+8)],data_in[`VWidth*(`APPRam_depth*28+9)-1:`VWidth*(`APPRam_depth*28+8)],data_in[`VWidth*(`APPRam_depth*27+9)-1:`VWidth*(`APPRam_depth*27+8)],data_in[`VWidth*(`APPRam_depth*26+9)-1:`VWidth*(`APPRam_depth*26+8)],data_in[`VWidth*(`APPRam_depth*25+9)-1:`VWidth*(`APPRam_depth*25+8)],data_in[`VWidth*(`APPRam_depth*24+9)-1:`VWidth*(`APPRam_depth*24+8)],data_in[`VWidth*(`APPRam_depth*23+9)-1:`VWidth*(`APPRam_depth*23+8)],data_in[`VWidth*(`APPRam_depth*22+9)-1:`VWidth*(`APPRam_depth*22+8)],data_in[`VWidth*(`APPRam_depth*21+9)-1:`VWidth*(`APPRam_depth*21+8)],data_in[`VWidth*(`APPRam_depth*20+9)-1:`VWidth*(`APPRam_depth*20+8)],data_in[`VWidth*(`APPRam_depth*19+9)-1:`VWidth*(`APPRam_depth*19+8)],data_in[`VWidth*(`APPRam_depth*18+9)-1:`VWidth*(`APPRam_depth*18+8)],data_in[`VWidth*(`APPRam_depth*17+9)-1:`VWidth*(`APPRam_depth*17+8)],data_in[`VWidth*(`APPRam_depth*16+9)-1:`VWidth*(`APPRam_depth*16+8)],data_in[`VWidth*(`APPRam_depth*15+9)-1:`VWidth*(`APPRam_depth*15+8)],data_in[`VWidth*(`APPRam_depth*14+9)-1:`VWidth*(`APPRam_depth*14+8)],data_in[`VWidth*(`APPRam_depth*13+9)-1:`VWidth*(`APPRam_depth*13+8)],data_in[`VWidth*(`APPRam_depth*12+9)-1:`VWidth*(`APPRam_depth*12+8)],data_in[`VWidth*(`APPRam_depth*11+9)-1:`VWidth*(`APPRam_depth*11+8)],data_in[`VWidth*(`APPRam_depth*10+9)-1:`VWidth*(`APPRam_depth*10+8)],data_in[`VWidth*(`APPRam_depth*9+9)-1:`VWidth*(`APPRam_depth*9+8)],data_in[`VWidth*(`APPRam_depth*8+9)-1:`VWidth*(`APPRam_depth*8+8)],data_in[`VWidth*(`APPRam_depth*7+9)-1:`VWidth*(`APPRam_depth*7+8)],data_in[`VWidth*(`APPRam_depth*6+9)-1:`VWidth*(`APPRam_depth*6+8)],data_in[`VWidth*(`APPRam_depth*5+9)-1:`VWidth*(`APPRam_depth*5+8)],data_in[`VWidth*(`APPRam_depth*4+9)-1:`VWidth*(`APPRam_depth*4+8)],data_in[`VWidth*(`APPRam_depth*3+9)-1:`VWidth*(`APPRam_depth*3+8)],data_in[`VWidth*(`APPRam_depth*2+9)-1:`VWidth*(`APPRam_depth*2+8)],data_in[`VWidth*(`APPRam_depth*1+9)-1:`VWidth*(`APPRam_depth*1+8)],data_in[`VWidth*(`APPRam_depth*0+9)-1:`VWidth*(`APPRam_depth*0+8)]};
			end
			9:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+10)-1:`VWidth*(`APPRam_depth*31+9)],data_in[`VWidth*(`APPRam_depth*30+10)-1:`VWidth*(`APPRam_depth*30+9)],data_in[`VWidth*(`APPRam_depth*29+10)-1:`VWidth*(`APPRam_depth*29+9)],data_in[`VWidth*(`APPRam_depth*28+10)-1:`VWidth*(`APPRam_depth*28+9)],data_in[`VWidth*(`APPRam_depth*27+10)-1:`VWidth*(`APPRam_depth*27+9)],data_in[`VWidth*(`APPRam_depth*26+10)-1:`VWidth*(`APPRam_depth*26+9)],data_in[`VWidth*(`APPRam_depth*25+10)-1:`VWidth*(`APPRam_depth*25+9)],data_in[`VWidth*(`APPRam_depth*24+10)-1:`VWidth*(`APPRam_depth*24+9)],data_in[`VWidth*(`APPRam_depth*23+10)-1:`VWidth*(`APPRam_depth*23+9)],data_in[`VWidth*(`APPRam_depth*22+10)-1:`VWidth*(`APPRam_depth*22+9)],data_in[`VWidth*(`APPRam_depth*21+10)-1:`VWidth*(`APPRam_depth*21+9)],data_in[`VWidth*(`APPRam_depth*20+10)-1:`VWidth*(`APPRam_depth*20+9)],data_in[`VWidth*(`APPRam_depth*19+10)-1:`VWidth*(`APPRam_depth*19+9)],data_in[`VWidth*(`APPRam_depth*18+10)-1:`VWidth*(`APPRam_depth*18+9)],data_in[`VWidth*(`APPRam_depth*17+10)-1:`VWidth*(`APPRam_depth*17+9)],data_in[`VWidth*(`APPRam_depth*16+10)-1:`VWidth*(`APPRam_depth*16+9)],data_in[`VWidth*(`APPRam_depth*15+10)-1:`VWidth*(`APPRam_depth*15+9)],data_in[`VWidth*(`APPRam_depth*14+10)-1:`VWidth*(`APPRam_depth*14+9)],data_in[`VWidth*(`APPRam_depth*13+10)-1:`VWidth*(`APPRam_depth*13+9)],data_in[`VWidth*(`APPRam_depth*12+10)-1:`VWidth*(`APPRam_depth*12+9)],data_in[`VWidth*(`APPRam_depth*11+10)-1:`VWidth*(`APPRam_depth*11+9)],data_in[`VWidth*(`APPRam_depth*10+10)-1:`VWidth*(`APPRam_depth*10+9)],data_in[`VWidth*(`APPRam_depth*9+10)-1:`VWidth*(`APPRam_depth*9+9)],data_in[`VWidth*(`APPRam_depth*8+10)-1:`VWidth*(`APPRam_depth*8+9)],data_in[`VWidth*(`APPRam_depth*7+10)-1:`VWidth*(`APPRam_depth*7+9)],data_in[`VWidth*(`APPRam_depth*6+10)-1:`VWidth*(`APPRam_depth*6+9)],data_in[`VWidth*(`APPRam_depth*5+10)-1:`VWidth*(`APPRam_depth*5+9)],data_in[`VWidth*(`APPRam_depth*4+10)-1:`VWidth*(`APPRam_depth*4+9)],data_in[`VWidth*(`APPRam_depth*3+10)-1:`VWidth*(`APPRam_depth*3+9)],data_in[`VWidth*(`APPRam_depth*2+10)-1:`VWidth*(`APPRam_depth*2+9)],data_in[`VWidth*(`APPRam_depth*1+10)-1:`VWidth*(`APPRam_depth*1+9)],data_in[`VWidth*(`APPRam_depth*0+10)-1:`VWidth*(`APPRam_depth*0+9)]};
			end
			10:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+11)-1:`VWidth*(`APPRam_depth*31+10)],data_in[`VWidth*(`APPRam_depth*30+11)-1:`VWidth*(`APPRam_depth*30+10)],data_in[`VWidth*(`APPRam_depth*29+11)-1:`VWidth*(`APPRam_depth*29+10)],data_in[`VWidth*(`APPRam_depth*28+11)-1:`VWidth*(`APPRam_depth*28+10)],data_in[`VWidth*(`APPRam_depth*27+11)-1:`VWidth*(`APPRam_depth*27+10)],data_in[`VWidth*(`APPRam_depth*26+11)-1:`VWidth*(`APPRam_depth*26+10)],data_in[`VWidth*(`APPRam_depth*25+11)-1:`VWidth*(`APPRam_depth*25+10)],data_in[`VWidth*(`APPRam_depth*24+11)-1:`VWidth*(`APPRam_depth*24+10)],data_in[`VWidth*(`APPRam_depth*23+11)-1:`VWidth*(`APPRam_depth*23+10)],data_in[`VWidth*(`APPRam_depth*22+11)-1:`VWidth*(`APPRam_depth*22+10)],data_in[`VWidth*(`APPRam_depth*21+11)-1:`VWidth*(`APPRam_depth*21+10)],data_in[`VWidth*(`APPRam_depth*20+11)-1:`VWidth*(`APPRam_depth*20+10)],data_in[`VWidth*(`APPRam_depth*19+11)-1:`VWidth*(`APPRam_depth*19+10)],data_in[`VWidth*(`APPRam_depth*18+11)-1:`VWidth*(`APPRam_depth*18+10)],data_in[`VWidth*(`APPRam_depth*17+11)-1:`VWidth*(`APPRam_depth*17+10)],data_in[`VWidth*(`APPRam_depth*16+11)-1:`VWidth*(`APPRam_depth*16+10)],data_in[`VWidth*(`APPRam_depth*15+11)-1:`VWidth*(`APPRam_depth*15+10)],data_in[`VWidth*(`APPRam_depth*14+11)-1:`VWidth*(`APPRam_depth*14+10)],data_in[`VWidth*(`APPRam_depth*13+11)-1:`VWidth*(`APPRam_depth*13+10)],data_in[`VWidth*(`APPRam_depth*12+11)-1:`VWidth*(`APPRam_depth*12+10)],data_in[`VWidth*(`APPRam_depth*11+11)-1:`VWidth*(`APPRam_depth*11+10)],data_in[`VWidth*(`APPRam_depth*10+11)-1:`VWidth*(`APPRam_depth*10+10)],data_in[`VWidth*(`APPRam_depth*9+11)-1:`VWidth*(`APPRam_depth*9+10)],data_in[`VWidth*(`APPRam_depth*8+11)-1:`VWidth*(`APPRam_depth*8+10)],data_in[`VWidth*(`APPRam_depth*7+11)-1:`VWidth*(`APPRam_depth*7+10)],data_in[`VWidth*(`APPRam_depth*6+11)-1:`VWidth*(`APPRam_depth*6+10)],data_in[`VWidth*(`APPRam_depth*5+11)-1:`VWidth*(`APPRam_depth*5+10)],data_in[`VWidth*(`APPRam_depth*4+11)-1:`VWidth*(`APPRam_depth*4+10)],data_in[`VWidth*(`APPRam_depth*3+11)-1:`VWidth*(`APPRam_depth*3+10)],data_in[`VWidth*(`APPRam_depth*2+11)-1:`VWidth*(`APPRam_depth*2+10)],data_in[`VWidth*(`APPRam_depth*1+11)-1:`VWidth*(`APPRam_depth*1+10)],data_in[`VWidth*(`APPRam_depth*0+11)-1:`VWidth*(`APPRam_depth*0+10)]};
			end
			11:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+12)-1:`VWidth*(`APPRam_depth*31+11)],data_in[`VWidth*(`APPRam_depth*30+12)-1:`VWidth*(`APPRam_depth*30+11)],data_in[`VWidth*(`APPRam_depth*29+12)-1:`VWidth*(`APPRam_depth*29+11)],data_in[`VWidth*(`APPRam_depth*28+12)-1:`VWidth*(`APPRam_depth*28+11)],data_in[`VWidth*(`APPRam_depth*27+12)-1:`VWidth*(`APPRam_depth*27+11)],data_in[`VWidth*(`APPRam_depth*26+12)-1:`VWidth*(`APPRam_depth*26+11)],data_in[`VWidth*(`APPRam_depth*25+12)-1:`VWidth*(`APPRam_depth*25+11)],data_in[`VWidth*(`APPRam_depth*24+12)-1:`VWidth*(`APPRam_depth*24+11)],data_in[`VWidth*(`APPRam_depth*23+12)-1:`VWidth*(`APPRam_depth*23+11)],data_in[`VWidth*(`APPRam_depth*22+12)-1:`VWidth*(`APPRam_depth*22+11)],data_in[`VWidth*(`APPRam_depth*21+12)-1:`VWidth*(`APPRam_depth*21+11)],data_in[`VWidth*(`APPRam_depth*20+12)-1:`VWidth*(`APPRam_depth*20+11)],data_in[`VWidth*(`APPRam_depth*19+12)-1:`VWidth*(`APPRam_depth*19+11)],data_in[`VWidth*(`APPRam_depth*18+12)-1:`VWidth*(`APPRam_depth*18+11)],data_in[`VWidth*(`APPRam_depth*17+12)-1:`VWidth*(`APPRam_depth*17+11)],data_in[`VWidth*(`APPRam_depth*16+12)-1:`VWidth*(`APPRam_depth*16+11)],data_in[`VWidth*(`APPRam_depth*15+12)-1:`VWidth*(`APPRam_depth*15+11)],data_in[`VWidth*(`APPRam_depth*14+12)-1:`VWidth*(`APPRam_depth*14+11)],data_in[`VWidth*(`APPRam_depth*13+12)-1:`VWidth*(`APPRam_depth*13+11)],data_in[`VWidth*(`APPRam_depth*12+12)-1:`VWidth*(`APPRam_depth*12+11)],data_in[`VWidth*(`APPRam_depth*11+12)-1:`VWidth*(`APPRam_depth*11+11)],data_in[`VWidth*(`APPRam_depth*10+12)-1:`VWidth*(`APPRam_depth*10+11)],data_in[`VWidth*(`APPRam_depth*9+12)-1:`VWidth*(`APPRam_depth*9+11)],data_in[`VWidth*(`APPRam_depth*8+12)-1:`VWidth*(`APPRam_depth*8+11)],data_in[`VWidth*(`APPRam_depth*7+12)-1:`VWidth*(`APPRam_depth*7+11)],data_in[`VWidth*(`APPRam_depth*6+12)-1:`VWidth*(`APPRam_depth*6+11)],data_in[`VWidth*(`APPRam_depth*5+12)-1:`VWidth*(`APPRam_depth*5+11)],data_in[`VWidth*(`APPRam_depth*4+12)-1:`VWidth*(`APPRam_depth*4+11)],data_in[`VWidth*(`APPRam_depth*3+12)-1:`VWidth*(`APPRam_depth*3+11)],data_in[`VWidth*(`APPRam_depth*2+12)-1:`VWidth*(`APPRam_depth*2+11)],data_in[`VWidth*(`APPRam_depth*1+12)-1:`VWidth*(`APPRam_depth*1+11)],data_in[`VWidth*(`APPRam_depth*0+12)-1:`VWidth*(`APPRam_depth*0+11)]};
			end
			12:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+13)-1:`VWidth*(`APPRam_depth*31+12)],data_in[`VWidth*(`APPRam_depth*30+13)-1:`VWidth*(`APPRam_depth*30+12)],data_in[`VWidth*(`APPRam_depth*29+13)-1:`VWidth*(`APPRam_depth*29+12)],data_in[`VWidth*(`APPRam_depth*28+13)-1:`VWidth*(`APPRam_depth*28+12)],data_in[`VWidth*(`APPRam_depth*27+13)-1:`VWidth*(`APPRam_depth*27+12)],data_in[`VWidth*(`APPRam_depth*26+13)-1:`VWidth*(`APPRam_depth*26+12)],data_in[`VWidth*(`APPRam_depth*25+13)-1:`VWidth*(`APPRam_depth*25+12)],data_in[`VWidth*(`APPRam_depth*24+13)-1:`VWidth*(`APPRam_depth*24+12)],data_in[`VWidth*(`APPRam_depth*23+13)-1:`VWidth*(`APPRam_depth*23+12)],data_in[`VWidth*(`APPRam_depth*22+13)-1:`VWidth*(`APPRam_depth*22+12)],data_in[`VWidth*(`APPRam_depth*21+13)-1:`VWidth*(`APPRam_depth*21+12)],data_in[`VWidth*(`APPRam_depth*20+13)-1:`VWidth*(`APPRam_depth*20+12)],data_in[`VWidth*(`APPRam_depth*19+13)-1:`VWidth*(`APPRam_depth*19+12)],data_in[`VWidth*(`APPRam_depth*18+13)-1:`VWidth*(`APPRam_depth*18+12)],data_in[`VWidth*(`APPRam_depth*17+13)-1:`VWidth*(`APPRam_depth*17+12)],data_in[`VWidth*(`APPRam_depth*16+13)-1:`VWidth*(`APPRam_depth*16+12)],data_in[`VWidth*(`APPRam_depth*15+13)-1:`VWidth*(`APPRam_depth*15+12)],data_in[`VWidth*(`APPRam_depth*14+13)-1:`VWidth*(`APPRam_depth*14+12)],data_in[`VWidth*(`APPRam_depth*13+13)-1:`VWidth*(`APPRam_depth*13+12)],data_in[`VWidth*(`APPRam_depth*12+13)-1:`VWidth*(`APPRam_depth*12+12)],data_in[`VWidth*(`APPRam_depth*11+13)-1:`VWidth*(`APPRam_depth*11+12)],data_in[`VWidth*(`APPRam_depth*10+13)-1:`VWidth*(`APPRam_depth*10+12)],data_in[`VWidth*(`APPRam_depth*9+13)-1:`VWidth*(`APPRam_depth*9+12)],data_in[`VWidth*(`APPRam_depth*8+13)-1:`VWidth*(`APPRam_depth*8+12)],data_in[`VWidth*(`APPRam_depth*7+13)-1:`VWidth*(`APPRam_depth*7+12)],data_in[`VWidth*(`APPRam_depth*6+13)-1:`VWidth*(`APPRam_depth*6+12)],data_in[`VWidth*(`APPRam_depth*5+13)-1:`VWidth*(`APPRam_depth*5+12)],data_in[`VWidth*(`APPRam_depth*4+13)-1:`VWidth*(`APPRam_depth*4+12)],data_in[`VWidth*(`APPRam_depth*3+13)-1:`VWidth*(`APPRam_depth*3+12)],data_in[`VWidth*(`APPRam_depth*2+13)-1:`VWidth*(`APPRam_depth*2+12)],data_in[`VWidth*(`APPRam_depth*1+13)-1:`VWidth*(`APPRam_depth*1+12)],data_in[`VWidth*(`APPRam_depth*0+13)-1:`VWidth*(`APPRam_depth*0+12)]};
			end
			13:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+14)-1:`VWidth*(`APPRam_depth*31+13)],data_in[`VWidth*(`APPRam_depth*30+14)-1:`VWidth*(`APPRam_depth*30+13)],data_in[`VWidth*(`APPRam_depth*29+14)-1:`VWidth*(`APPRam_depth*29+13)],data_in[`VWidth*(`APPRam_depth*28+14)-1:`VWidth*(`APPRam_depth*28+13)],data_in[`VWidth*(`APPRam_depth*27+14)-1:`VWidth*(`APPRam_depth*27+13)],data_in[`VWidth*(`APPRam_depth*26+14)-1:`VWidth*(`APPRam_depth*26+13)],data_in[`VWidth*(`APPRam_depth*25+14)-1:`VWidth*(`APPRam_depth*25+13)],data_in[`VWidth*(`APPRam_depth*24+14)-1:`VWidth*(`APPRam_depth*24+13)],data_in[`VWidth*(`APPRam_depth*23+14)-1:`VWidth*(`APPRam_depth*23+13)],data_in[`VWidth*(`APPRam_depth*22+14)-1:`VWidth*(`APPRam_depth*22+13)],data_in[`VWidth*(`APPRam_depth*21+14)-1:`VWidth*(`APPRam_depth*21+13)],data_in[`VWidth*(`APPRam_depth*20+14)-1:`VWidth*(`APPRam_depth*20+13)],data_in[`VWidth*(`APPRam_depth*19+14)-1:`VWidth*(`APPRam_depth*19+13)],data_in[`VWidth*(`APPRam_depth*18+14)-1:`VWidth*(`APPRam_depth*18+13)],data_in[`VWidth*(`APPRam_depth*17+14)-1:`VWidth*(`APPRam_depth*17+13)],data_in[`VWidth*(`APPRam_depth*16+14)-1:`VWidth*(`APPRam_depth*16+13)],data_in[`VWidth*(`APPRam_depth*15+14)-1:`VWidth*(`APPRam_depth*15+13)],data_in[`VWidth*(`APPRam_depth*14+14)-1:`VWidth*(`APPRam_depth*14+13)],data_in[`VWidth*(`APPRam_depth*13+14)-1:`VWidth*(`APPRam_depth*13+13)],data_in[`VWidth*(`APPRam_depth*12+14)-1:`VWidth*(`APPRam_depth*12+13)],data_in[`VWidth*(`APPRam_depth*11+14)-1:`VWidth*(`APPRam_depth*11+13)],data_in[`VWidth*(`APPRam_depth*10+14)-1:`VWidth*(`APPRam_depth*10+13)],data_in[`VWidth*(`APPRam_depth*9+14)-1:`VWidth*(`APPRam_depth*9+13)],data_in[`VWidth*(`APPRam_depth*8+14)-1:`VWidth*(`APPRam_depth*8+13)],data_in[`VWidth*(`APPRam_depth*7+14)-1:`VWidth*(`APPRam_depth*7+13)],data_in[`VWidth*(`APPRam_depth*6+14)-1:`VWidth*(`APPRam_depth*6+13)],data_in[`VWidth*(`APPRam_depth*5+14)-1:`VWidth*(`APPRam_depth*5+13)],data_in[`VWidth*(`APPRam_depth*4+14)-1:`VWidth*(`APPRam_depth*4+13)],data_in[`VWidth*(`APPRam_depth*3+14)-1:`VWidth*(`APPRam_depth*3+13)],data_in[`VWidth*(`APPRam_depth*2+14)-1:`VWidth*(`APPRam_depth*2+13)],data_in[`VWidth*(`APPRam_depth*1+14)-1:`VWidth*(`APPRam_depth*1+13)],data_in[`VWidth*(`APPRam_depth*0+14)-1:`VWidth*(`APPRam_depth*0+13)]};
			end
			14:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+15)-1:`VWidth*(`APPRam_depth*31+14)],data_in[`VWidth*(`APPRam_depth*30+15)-1:`VWidth*(`APPRam_depth*30+14)],data_in[`VWidth*(`APPRam_depth*29+15)-1:`VWidth*(`APPRam_depth*29+14)],data_in[`VWidth*(`APPRam_depth*28+15)-1:`VWidth*(`APPRam_depth*28+14)],data_in[`VWidth*(`APPRam_depth*27+15)-1:`VWidth*(`APPRam_depth*27+14)],data_in[`VWidth*(`APPRam_depth*26+15)-1:`VWidth*(`APPRam_depth*26+14)],data_in[`VWidth*(`APPRam_depth*25+15)-1:`VWidth*(`APPRam_depth*25+14)],data_in[`VWidth*(`APPRam_depth*24+15)-1:`VWidth*(`APPRam_depth*24+14)],data_in[`VWidth*(`APPRam_depth*23+15)-1:`VWidth*(`APPRam_depth*23+14)],data_in[`VWidth*(`APPRam_depth*22+15)-1:`VWidth*(`APPRam_depth*22+14)],data_in[`VWidth*(`APPRam_depth*21+15)-1:`VWidth*(`APPRam_depth*21+14)],data_in[`VWidth*(`APPRam_depth*20+15)-1:`VWidth*(`APPRam_depth*20+14)],data_in[`VWidth*(`APPRam_depth*19+15)-1:`VWidth*(`APPRam_depth*19+14)],data_in[`VWidth*(`APPRam_depth*18+15)-1:`VWidth*(`APPRam_depth*18+14)],data_in[`VWidth*(`APPRam_depth*17+15)-1:`VWidth*(`APPRam_depth*17+14)],data_in[`VWidth*(`APPRam_depth*16+15)-1:`VWidth*(`APPRam_depth*16+14)],data_in[`VWidth*(`APPRam_depth*15+15)-1:`VWidth*(`APPRam_depth*15+14)],data_in[`VWidth*(`APPRam_depth*14+15)-1:`VWidth*(`APPRam_depth*14+14)],data_in[`VWidth*(`APPRam_depth*13+15)-1:`VWidth*(`APPRam_depth*13+14)],data_in[`VWidth*(`APPRam_depth*12+15)-1:`VWidth*(`APPRam_depth*12+14)],data_in[`VWidth*(`APPRam_depth*11+15)-1:`VWidth*(`APPRam_depth*11+14)],data_in[`VWidth*(`APPRam_depth*10+15)-1:`VWidth*(`APPRam_depth*10+14)],data_in[`VWidth*(`APPRam_depth*9+15)-1:`VWidth*(`APPRam_depth*9+14)],data_in[`VWidth*(`APPRam_depth*8+15)-1:`VWidth*(`APPRam_depth*8+14)],data_in[`VWidth*(`APPRam_depth*7+15)-1:`VWidth*(`APPRam_depth*7+14)],data_in[`VWidth*(`APPRam_depth*6+15)-1:`VWidth*(`APPRam_depth*6+14)],data_in[`VWidth*(`APPRam_depth*5+15)-1:`VWidth*(`APPRam_depth*5+14)],data_in[`VWidth*(`APPRam_depth*4+15)-1:`VWidth*(`APPRam_depth*4+14)],data_in[`VWidth*(`APPRam_depth*3+15)-1:`VWidth*(`APPRam_depth*3+14)],data_in[`VWidth*(`APPRam_depth*2+15)-1:`VWidth*(`APPRam_depth*2+14)],data_in[`VWidth*(`APPRam_depth*1+15)-1:`VWidth*(`APPRam_depth*1+14)],data_in[`VWidth*(`APPRam_depth*0+15)-1:`VWidth*(`APPRam_depth*0+14)]};
			end
			15:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+16)-1:`VWidth*(`APPRam_depth*31+15)],data_in[`VWidth*(`APPRam_depth*30+16)-1:`VWidth*(`APPRam_depth*30+15)],data_in[`VWidth*(`APPRam_depth*29+16)-1:`VWidth*(`APPRam_depth*29+15)],data_in[`VWidth*(`APPRam_depth*28+16)-1:`VWidth*(`APPRam_depth*28+15)],data_in[`VWidth*(`APPRam_depth*27+16)-1:`VWidth*(`APPRam_depth*27+15)],data_in[`VWidth*(`APPRam_depth*26+16)-1:`VWidth*(`APPRam_depth*26+15)],data_in[`VWidth*(`APPRam_depth*25+16)-1:`VWidth*(`APPRam_depth*25+15)],data_in[`VWidth*(`APPRam_depth*24+16)-1:`VWidth*(`APPRam_depth*24+15)],data_in[`VWidth*(`APPRam_depth*23+16)-1:`VWidth*(`APPRam_depth*23+15)],data_in[`VWidth*(`APPRam_depth*22+16)-1:`VWidth*(`APPRam_depth*22+15)],data_in[`VWidth*(`APPRam_depth*21+16)-1:`VWidth*(`APPRam_depth*21+15)],data_in[`VWidth*(`APPRam_depth*20+16)-1:`VWidth*(`APPRam_depth*20+15)],data_in[`VWidth*(`APPRam_depth*19+16)-1:`VWidth*(`APPRam_depth*19+15)],data_in[`VWidth*(`APPRam_depth*18+16)-1:`VWidth*(`APPRam_depth*18+15)],data_in[`VWidth*(`APPRam_depth*17+16)-1:`VWidth*(`APPRam_depth*17+15)],data_in[`VWidth*(`APPRam_depth*16+16)-1:`VWidth*(`APPRam_depth*16+15)],data_in[`VWidth*(`APPRam_depth*15+16)-1:`VWidth*(`APPRam_depth*15+15)],data_in[`VWidth*(`APPRam_depth*14+16)-1:`VWidth*(`APPRam_depth*14+15)],data_in[`VWidth*(`APPRam_depth*13+16)-1:`VWidth*(`APPRam_depth*13+15)],data_in[`VWidth*(`APPRam_depth*12+16)-1:`VWidth*(`APPRam_depth*12+15)],data_in[`VWidth*(`APPRam_depth*11+16)-1:`VWidth*(`APPRam_depth*11+15)],data_in[`VWidth*(`APPRam_depth*10+16)-1:`VWidth*(`APPRam_depth*10+15)],data_in[`VWidth*(`APPRam_depth*9+16)-1:`VWidth*(`APPRam_depth*9+15)],data_in[`VWidth*(`APPRam_depth*8+16)-1:`VWidth*(`APPRam_depth*8+15)],data_in[`VWidth*(`APPRam_depth*7+16)-1:`VWidth*(`APPRam_depth*7+15)],data_in[`VWidth*(`APPRam_depth*6+16)-1:`VWidth*(`APPRam_depth*6+15)],data_in[`VWidth*(`APPRam_depth*5+16)-1:`VWidth*(`APPRam_depth*5+15)],data_in[`VWidth*(`APPRam_depth*4+16)-1:`VWidth*(`APPRam_depth*4+15)],data_in[`VWidth*(`APPRam_depth*3+16)-1:`VWidth*(`APPRam_depth*3+15)],data_in[`VWidth*(`APPRam_depth*2+16)-1:`VWidth*(`APPRam_depth*2+15)],data_in[`VWidth*(`APPRam_depth*1+16)-1:`VWidth*(`APPRam_depth*1+15)],data_in[`VWidth*(`APPRam_depth*0+16)-1:`VWidth*(`APPRam_depth*0+15)]};
			end

			default:
			begin
				data_out <= 0;
			end
		endcase
	end
	else
	begin
		data_out <= 0;
	end
end


endmodule