`include "Decoder_Parameters.v"
module get_msgini(
    input clk,
    input rst_n,
    input [`Zc*`VWidth-1:0] data_in, //输入目的是分割一个方阵的元素为Zc/DPU_num组
    input [`APP_addr_width-2:0] addr_in,
	input en_in,
    output reg [`inNum*`VWidth-1:0] data_out //输出32长度，就是DPU并行度的长度
	// output reg [`APP_addr_width-2:0] addr_out
);

reg [`APP_addr_width-2:0] addr_in_D0;
// always @(posedge clk or negedge rst_n)
// begin
// 	if(!rst_n)
// 	begin
// 		addr_out <= 0;
// 	end
// 	else
// 	begin
// 		addr_out <= addr_in;
// 	end
// end

always @(posedge clk or negedge rst_n)
begin
	if(!rst_n)
	begin
		addr_in_D0 <= 0;
	end
	else
	begin
		addr_in_D0 <= addr_in;
	end
end

always @(posedge clk or negedge rst_n)
begin
	if(!rst_n)
	begin
		data_out <= 0;
	end
	else if(en_in)
	begin
		case(addr_in)
			0:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+1)-1:`VWidth*(`APPRam_depth*31+0)],data_in[`VWidth*(`APPRam_depth*30+1)-1:`VWidth*(`APPRam_depth*30+0)],data_in[`VWidth*(`APPRam_depth*29+1)-1:`VWidth*(`APPRam_depth*29+0)],data_in[`VWidth*(`APPRam_depth*28+1)-1:`VWidth*(`APPRam_depth*28+0)],data_in[`VWidth*(`APPRam_depth*27+1)-1:`VWidth*(`APPRam_depth*27+0)],data_in[`VWidth*(`APPRam_depth*26+1)-1:`VWidth*(`APPRam_depth*26+0)],data_in[`VWidth*(`APPRam_depth*25+1)-1:`VWidth*(`APPRam_depth*25+0)],data_in[`VWidth*(`APPRam_depth*24+1)-1:`VWidth*(`APPRam_depth*24+0)],data_in[`VWidth*(`APPRam_depth*23+1)-1:`VWidth*(`APPRam_depth*23+0)],data_in[`VWidth*(`APPRam_depth*22+1)-1:`VWidth*(`APPRam_depth*22+0)],data_in[`VWidth*(`APPRam_depth*21+1)-1:`VWidth*(`APPRam_depth*21+0)],data_in[`VWidth*(`APPRam_depth*20+1)-1:`VWidth*(`APPRam_depth*20+0)],data_in[`VWidth*(`APPRam_depth*19+1)-1:`VWidth*(`APPRam_depth*19+0)],data_in[`VWidth*(`APPRam_depth*18+1)-1:`VWidth*(`APPRam_depth*18+0)],data_in[`VWidth*(`APPRam_depth*17+1)-1:`VWidth*(`APPRam_depth*17+0)],data_in[`VWidth*(`APPRam_depth*16+1)-1:`VWidth*(`APPRam_depth*16+0)],data_in[`VWidth*(`APPRam_depth*15+1)-1:`VWidth*(`APPRam_depth*15+0)],data_in[`VWidth*(`APPRam_depth*14+1)-1:`VWidth*(`APPRam_depth*14+0)],data_in[`VWidth*(`APPRam_depth*13+1)-1:`VWidth*(`APPRam_depth*13+0)],data_in[`VWidth*(`APPRam_depth*12+1)-1:`VWidth*(`APPRam_depth*12+0)],data_in[`VWidth*(`APPRam_depth*11+1)-1:`VWidth*(`APPRam_depth*11+0)],data_in[`VWidth*(`APPRam_depth*10+1)-1:`VWidth*(`APPRam_depth*10+0)],data_in[`VWidth*(`APPRam_depth*9+1)-1:`VWidth*(`APPRam_depth*9+0)],data_in[`VWidth*(`APPRam_depth*8+1)-1:`VWidth*(`APPRam_depth*8+0)],data_in[`VWidth*(`APPRam_depth*7+1)-1:`VWidth*(`APPRam_depth*7+0)],data_in[`VWidth*(`APPRam_depth*6+1)-1:`VWidth*(`APPRam_depth*6+0)],data_in[`VWidth*(`APPRam_depth*5+1)-1:`VWidth*(`APPRam_depth*5+0)],data_in[`VWidth*(`APPRam_depth*4+1)-1:`VWidth*(`APPRam_depth*4+0)],data_in[`VWidth*(`APPRam_depth*3+1)-1:`VWidth*(`APPRam_depth*3+0)],data_in[`VWidth*(`APPRam_depth*2+1)-1:`VWidth*(`APPRam_depth*2+0)],data_in[`VWidth*(`APPRam_depth*1+1)-1:`VWidth*(`APPRam_depth*1+0)],data_in[`VWidth*(`APPRam_depth*0+1)-1:`VWidth*(`APPRam_depth*0+0)]};
			end
			1:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+2)-1:`VWidth*(`APPRam_depth*31+1)],data_in[`VWidth*(`APPRam_depth*30+2)-1:`VWidth*(`APPRam_depth*30+1)],data_in[`VWidth*(`APPRam_depth*29+2)-1:`VWidth*(`APPRam_depth*29+1)],data_in[`VWidth*(`APPRam_depth*28+2)-1:`VWidth*(`APPRam_depth*28+1)],data_in[`VWidth*(`APPRam_depth*27+2)-1:`VWidth*(`APPRam_depth*27+1)],data_in[`VWidth*(`APPRam_depth*26+2)-1:`VWidth*(`APPRam_depth*26+1)],data_in[`VWidth*(`APPRam_depth*25+2)-1:`VWidth*(`APPRam_depth*25+1)],data_in[`VWidth*(`APPRam_depth*24+2)-1:`VWidth*(`APPRam_depth*24+1)],data_in[`VWidth*(`APPRam_depth*23+2)-1:`VWidth*(`APPRam_depth*23+1)],data_in[`VWidth*(`APPRam_depth*22+2)-1:`VWidth*(`APPRam_depth*22+1)],data_in[`VWidth*(`APPRam_depth*21+2)-1:`VWidth*(`APPRam_depth*21+1)],data_in[`VWidth*(`APPRam_depth*20+2)-1:`VWidth*(`APPRam_depth*20+1)],data_in[`VWidth*(`APPRam_depth*19+2)-1:`VWidth*(`APPRam_depth*19+1)],data_in[`VWidth*(`APPRam_depth*18+2)-1:`VWidth*(`APPRam_depth*18+1)],data_in[`VWidth*(`APPRam_depth*17+2)-1:`VWidth*(`APPRam_depth*17+1)],data_in[`VWidth*(`APPRam_depth*16+2)-1:`VWidth*(`APPRam_depth*16+1)],data_in[`VWidth*(`APPRam_depth*15+2)-1:`VWidth*(`APPRam_depth*15+1)],data_in[`VWidth*(`APPRam_depth*14+2)-1:`VWidth*(`APPRam_depth*14+1)],data_in[`VWidth*(`APPRam_depth*13+2)-1:`VWidth*(`APPRam_depth*13+1)],data_in[`VWidth*(`APPRam_depth*12+2)-1:`VWidth*(`APPRam_depth*12+1)],data_in[`VWidth*(`APPRam_depth*11+2)-1:`VWidth*(`APPRam_depth*11+1)],data_in[`VWidth*(`APPRam_depth*10+2)-1:`VWidth*(`APPRam_depth*10+1)],data_in[`VWidth*(`APPRam_depth*9+2)-1:`VWidth*(`APPRam_depth*9+1)],data_in[`VWidth*(`APPRam_depth*8+2)-1:`VWidth*(`APPRam_depth*8+1)],data_in[`VWidth*(`APPRam_depth*7+2)-1:`VWidth*(`APPRam_depth*7+1)],data_in[`VWidth*(`APPRam_depth*6+2)-1:`VWidth*(`APPRam_depth*6+1)],data_in[`VWidth*(`APPRam_depth*5+2)-1:`VWidth*(`APPRam_depth*5+1)],data_in[`VWidth*(`APPRam_depth*4+2)-1:`VWidth*(`APPRam_depth*4+1)],data_in[`VWidth*(`APPRam_depth*3+2)-1:`VWidth*(`APPRam_depth*3+1)],data_in[`VWidth*(`APPRam_depth*2+2)-1:`VWidth*(`APPRam_depth*2+1)],data_in[`VWidth*(`APPRam_depth*1+2)-1:`VWidth*(`APPRam_depth*1+1)],data_in[`VWidth*(`APPRam_depth*0+2)-1:`VWidth*(`APPRam_depth*0+1)]};
			end
			2:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+3)-1:`VWidth*(`APPRam_depth*31+2)],data_in[`VWidth*(`APPRam_depth*30+3)-1:`VWidth*(`APPRam_depth*30+2)],data_in[`VWidth*(`APPRam_depth*29+3)-1:`VWidth*(`APPRam_depth*29+2)],data_in[`VWidth*(`APPRam_depth*28+3)-1:`VWidth*(`APPRam_depth*28+2)],data_in[`VWidth*(`APPRam_depth*27+3)-1:`VWidth*(`APPRam_depth*27+2)],data_in[`VWidth*(`APPRam_depth*26+3)-1:`VWidth*(`APPRam_depth*26+2)],data_in[`VWidth*(`APPRam_depth*25+3)-1:`VWidth*(`APPRam_depth*25+2)],data_in[`VWidth*(`APPRam_depth*24+3)-1:`VWidth*(`APPRam_depth*24+2)],data_in[`VWidth*(`APPRam_depth*23+3)-1:`VWidth*(`APPRam_depth*23+2)],data_in[`VWidth*(`APPRam_depth*22+3)-1:`VWidth*(`APPRam_depth*22+2)],data_in[`VWidth*(`APPRam_depth*21+3)-1:`VWidth*(`APPRam_depth*21+2)],data_in[`VWidth*(`APPRam_depth*20+3)-1:`VWidth*(`APPRam_depth*20+2)],data_in[`VWidth*(`APPRam_depth*19+3)-1:`VWidth*(`APPRam_depth*19+2)],data_in[`VWidth*(`APPRam_depth*18+3)-1:`VWidth*(`APPRam_depth*18+2)],data_in[`VWidth*(`APPRam_depth*17+3)-1:`VWidth*(`APPRam_depth*17+2)],data_in[`VWidth*(`APPRam_depth*16+3)-1:`VWidth*(`APPRam_depth*16+2)],data_in[`VWidth*(`APPRam_depth*15+3)-1:`VWidth*(`APPRam_depth*15+2)],data_in[`VWidth*(`APPRam_depth*14+3)-1:`VWidth*(`APPRam_depth*14+2)],data_in[`VWidth*(`APPRam_depth*13+3)-1:`VWidth*(`APPRam_depth*13+2)],data_in[`VWidth*(`APPRam_depth*12+3)-1:`VWidth*(`APPRam_depth*12+2)],data_in[`VWidth*(`APPRam_depth*11+3)-1:`VWidth*(`APPRam_depth*11+2)],data_in[`VWidth*(`APPRam_depth*10+3)-1:`VWidth*(`APPRam_depth*10+2)],data_in[`VWidth*(`APPRam_depth*9+3)-1:`VWidth*(`APPRam_depth*9+2)],data_in[`VWidth*(`APPRam_depth*8+3)-1:`VWidth*(`APPRam_depth*8+2)],data_in[`VWidth*(`APPRam_depth*7+3)-1:`VWidth*(`APPRam_depth*7+2)],data_in[`VWidth*(`APPRam_depth*6+3)-1:`VWidth*(`APPRam_depth*6+2)],data_in[`VWidth*(`APPRam_depth*5+3)-1:`VWidth*(`APPRam_depth*5+2)],data_in[`VWidth*(`APPRam_depth*4+3)-1:`VWidth*(`APPRam_depth*4+2)],data_in[`VWidth*(`APPRam_depth*3+3)-1:`VWidth*(`APPRam_depth*3+2)],data_in[`VWidth*(`APPRam_depth*2+3)-1:`VWidth*(`APPRam_depth*2+2)],data_in[`VWidth*(`APPRam_depth*1+3)-1:`VWidth*(`APPRam_depth*1+2)],data_in[`VWidth*(`APPRam_depth*0+3)-1:`VWidth*(`APPRam_depth*0+2)]};
			end
			3:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+4)-1:`VWidth*(`APPRam_depth*31+3)],data_in[`VWidth*(`APPRam_depth*30+4)-1:`VWidth*(`APPRam_depth*30+3)],data_in[`VWidth*(`APPRam_depth*29+4)-1:`VWidth*(`APPRam_depth*29+3)],data_in[`VWidth*(`APPRam_depth*28+4)-1:`VWidth*(`APPRam_depth*28+3)],data_in[`VWidth*(`APPRam_depth*27+4)-1:`VWidth*(`APPRam_depth*27+3)],data_in[`VWidth*(`APPRam_depth*26+4)-1:`VWidth*(`APPRam_depth*26+3)],data_in[`VWidth*(`APPRam_depth*25+4)-1:`VWidth*(`APPRam_depth*25+3)],data_in[`VWidth*(`APPRam_depth*24+4)-1:`VWidth*(`APPRam_depth*24+3)],data_in[`VWidth*(`APPRam_depth*23+4)-1:`VWidth*(`APPRam_depth*23+3)],data_in[`VWidth*(`APPRam_depth*22+4)-1:`VWidth*(`APPRam_depth*22+3)],data_in[`VWidth*(`APPRam_depth*21+4)-1:`VWidth*(`APPRam_depth*21+3)],data_in[`VWidth*(`APPRam_depth*20+4)-1:`VWidth*(`APPRam_depth*20+3)],data_in[`VWidth*(`APPRam_depth*19+4)-1:`VWidth*(`APPRam_depth*19+3)],data_in[`VWidth*(`APPRam_depth*18+4)-1:`VWidth*(`APPRam_depth*18+3)],data_in[`VWidth*(`APPRam_depth*17+4)-1:`VWidth*(`APPRam_depth*17+3)],data_in[`VWidth*(`APPRam_depth*16+4)-1:`VWidth*(`APPRam_depth*16+3)],data_in[`VWidth*(`APPRam_depth*15+4)-1:`VWidth*(`APPRam_depth*15+3)],data_in[`VWidth*(`APPRam_depth*14+4)-1:`VWidth*(`APPRam_depth*14+3)],data_in[`VWidth*(`APPRam_depth*13+4)-1:`VWidth*(`APPRam_depth*13+3)],data_in[`VWidth*(`APPRam_depth*12+4)-1:`VWidth*(`APPRam_depth*12+3)],data_in[`VWidth*(`APPRam_depth*11+4)-1:`VWidth*(`APPRam_depth*11+3)],data_in[`VWidth*(`APPRam_depth*10+4)-1:`VWidth*(`APPRam_depth*10+3)],data_in[`VWidth*(`APPRam_depth*9+4)-1:`VWidth*(`APPRam_depth*9+3)],data_in[`VWidth*(`APPRam_depth*8+4)-1:`VWidth*(`APPRam_depth*8+3)],data_in[`VWidth*(`APPRam_depth*7+4)-1:`VWidth*(`APPRam_depth*7+3)],data_in[`VWidth*(`APPRam_depth*6+4)-1:`VWidth*(`APPRam_depth*6+3)],data_in[`VWidth*(`APPRam_depth*5+4)-1:`VWidth*(`APPRam_depth*5+3)],data_in[`VWidth*(`APPRam_depth*4+4)-1:`VWidth*(`APPRam_depth*4+3)],data_in[`VWidth*(`APPRam_depth*3+4)-1:`VWidth*(`APPRam_depth*3+3)],data_in[`VWidth*(`APPRam_depth*2+4)-1:`VWidth*(`APPRam_depth*2+3)],data_in[`VWidth*(`APPRam_depth*1+4)-1:`VWidth*(`APPRam_depth*1+3)],data_in[`VWidth*(`APPRam_depth*0+4)-1:`VWidth*(`APPRam_depth*0+3)]};
			end
			4:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+5)-1:`VWidth*(`APPRam_depth*31+4)],data_in[`VWidth*(`APPRam_depth*30+5)-1:`VWidth*(`APPRam_depth*30+4)],data_in[`VWidth*(`APPRam_depth*29+5)-1:`VWidth*(`APPRam_depth*29+4)],data_in[`VWidth*(`APPRam_depth*28+5)-1:`VWidth*(`APPRam_depth*28+4)],data_in[`VWidth*(`APPRam_depth*27+5)-1:`VWidth*(`APPRam_depth*27+4)],data_in[`VWidth*(`APPRam_depth*26+5)-1:`VWidth*(`APPRam_depth*26+4)],data_in[`VWidth*(`APPRam_depth*25+5)-1:`VWidth*(`APPRam_depth*25+4)],data_in[`VWidth*(`APPRam_depth*24+5)-1:`VWidth*(`APPRam_depth*24+4)],data_in[`VWidth*(`APPRam_depth*23+5)-1:`VWidth*(`APPRam_depth*23+4)],data_in[`VWidth*(`APPRam_depth*22+5)-1:`VWidth*(`APPRam_depth*22+4)],data_in[`VWidth*(`APPRam_depth*21+5)-1:`VWidth*(`APPRam_depth*21+4)],data_in[`VWidth*(`APPRam_depth*20+5)-1:`VWidth*(`APPRam_depth*20+4)],data_in[`VWidth*(`APPRam_depth*19+5)-1:`VWidth*(`APPRam_depth*19+4)],data_in[`VWidth*(`APPRam_depth*18+5)-1:`VWidth*(`APPRam_depth*18+4)],data_in[`VWidth*(`APPRam_depth*17+5)-1:`VWidth*(`APPRam_depth*17+4)],data_in[`VWidth*(`APPRam_depth*16+5)-1:`VWidth*(`APPRam_depth*16+4)],data_in[`VWidth*(`APPRam_depth*15+5)-1:`VWidth*(`APPRam_depth*15+4)],data_in[`VWidth*(`APPRam_depth*14+5)-1:`VWidth*(`APPRam_depth*14+4)],data_in[`VWidth*(`APPRam_depth*13+5)-1:`VWidth*(`APPRam_depth*13+4)],data_in[`VWidth*(`APPRam_depth*12+5)-1:`VWidth*(`APPRam_depth*12+4)],data_in[`VWidth*(`APPRam_depth*11+5)-1:`VWidth*(`APPRam_depth*11+4)],data_in[`VWidth*(`APPRam_depth*10+5)-1:`VWidth*(`APPRam_depth*10+4)],data_in[`VWidth*(`APPRam_depth*9+5)-1:`VWidth*(`APPRam_depth*9+4)],data_in[`VWidth*(`APPRam_depth*8+5)-1:`VWidth*(`APPRam_depth*8+4)],data_in[`VWidth*(`APPRam_depth*7+5)-1:`VWidth*(`APPRam_depth*7+4)],data_in[`VWidth*(`APPRam_depth*6+5)-1:`VWidth*(`APPRam_depth*6+4)],data_in[`VWidth*(`APPRam_depth*5+5)-1:`VWidth*(`APPRam_depth*5+4)],data_in[`VWidth*(`APPRam_depth*4+5)-1:`VWidth*(`APPRam_depth*4+4)],data_in[`VWidth*(`APPRam_depth*3+5)-1:`VWidth*(`APPRam_depth*3+4)],data_in[`VWidth*(`APPRam_depth*2+5)-1:`VWidth*(`APPRam_depth*2+4)],data_in[`VWidth*(`APPRam_depth*1+5)-1:`VWidth*(`APPRam_depth*1+4)],data_in[`VWidth*(`APPRam_depth*0+5)-1:`VWidth*(`APPRam_depth*0+4)]};
			end
			5:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+6)-1:`VWidth*(`APPRam_depth*31+5)],data_in[`VWidth*(`APPRam_depth*30+6)-1:`VWidth*(`APPRam_depth*30+5)],data_in[`VWidth*(`APPRam_depth*29+6)-1:`VWidth*(`APPRam_depth*29+5)],data_in[`VWidth*(`APPRam_depth*28+6)-1:`VWidth*(`APPRam_depth*28+5)],data_in[`VWidth*(`APPRam_depth*27+6)-1:`VWidth*(`APPRam_depth*27+5)],data_in[`VWidth*(`APPRam_depth*26+6)-1:`VWidth*(`APPRam_depth*26+5)],data_in[`VWidth*(`APPRam_depth*25+6)-1:`VWidth*(`APPRam_depth*25+5)],data_in[`VWidth*(`APPRam_depth*24+6)-1:`VWidth*(`APPRam_depth*24+5)],data_in[`VWidth*(`APPRam_depth*23+6)-1:`VWidth*(`APPRam_depth*23+5)],data_in[`VWidth*(`APPRam_depth*22+6)-1:`VWidth*(`APPRam_depth*22+5)],data_in[`VWidth*(`APPRam_depth*21+6)-1:`VWidth*(`APPRam_depth*21+5)],data_in[`VWidth*(`APPRam_depth*20+6)-1:`VWidth*(`APPRam_depth*20+5)],data_in[`VWidth*(`APPRam_depth*19+6)-1:`VWidth*(`APPRam_depth*19+5)],data_in[`VWidth*(`APPRam_depth*18+6)-1:`VWidth*(`APPRam_depth*18+5)],data_in[`VWidth*(`APPRam_depth*17+6)-1:`VWidth*(`APPRam_depth*17+5)],data_in[`VWidth*(`APPRam_depth*16+6)-1:`VWidth*(`APPRam_depth*16+5)],data_in[`VWidth*(`APPRam_depth*15+6)-1:`VWidth*(`APPRam_depth*15+5)],data_in[`VWidth*(`APPRam_depth*14+6)-1:`VWidth*(`APPRam_depth*14+5)],data_in[`VWidth*(`APPRam_depth*13+6)-1:`VWidth*(`APPRam_depth*13+5)],data_in[`VWidth*(`APPRam_depth*12+6)-1:`VWidth*(`APPRam_depth*12+5)],data_in[`VWidth*(`APPRam_depth*11+6)-1:`VWidth*(`APPRam_depth*11+5)],data_in[`VWidth*(`APPRam_depth*10+6)-1:`VWidth*(`APPRam_depth*10+5)],data_in[`VWidth*(`APPRam_depth*9+6)-1:`VWidth*(`APPRam_depth*9+5)],data_in[`VWidth*(`APPRam_depth*8+6)-1:`VWidth*(`APPRam_depth*8+5)],data_in[`VWidth*(`APPRam_depth*7+6)-1:`VWidth*(`APPRam_depth*7+5)],data_in[`VWidth*(`APPRam_depth*6+6)-1:`VWidth*(`APPRam_depth*6+5)],data_in[`VWidth*(`APPRam_depth*5+6)-1:`VWidth*(`APPRam_depth*5+5)],data_in[`VWidth*(`APPRam_depth*4+6)-1:`VWidth*(`APPRam_depth*4+5)],data_in[`VWidth*(`APPRam_depth*3+6)-1:`VWidth*(`APPRam_depth*3+5)],data_in[`VWidth*(`APPRam_depth*2+6)-1:`VWidth*(`APPRam_depth*2+5)],data_in[`VWidth*(`APPRam_depth*1+6)-1:`VWidth*(`APPRam_depth*1+5)],data_in[`VWidth*(`APPRam_depth*0+6)-1:`VWidth*(`APPRam_depth*0+5)]};
			end
			6:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+7)-1:`VWidth*(`APPRam_depth*31+6)],data_in[`VWidth*(`APPRam_depth*30+7)-1:`VWidth*(`APPRam_depth*30+6)],data_in[`VWidth*(`APPRam_depth*29+7)-1:`VWidth*(`APPRam_depth*29+6)],data_in[`VWidth*(`APPRam_depth*28+7)-1:`VWidth*(`APPRam_depth*28+6)],data_in[`VWidth*(`APPRam_depth*27+7)-1:`VWidth*(`APPRam_depth*27+6)],data_in[`VWidth*(`APPRam_depth*26+7)-1:`VWidth*(`APPRam_depth*26+6)],data_in[`VWidth*(`APPRam_depth*25+7)-1:`VWidth*(`APPRam_depth*25+6)],data_in[`VWidth*(`APPRam_depth*24+7)-1:`VWidth*(`APPRam_depth*24+6)],data_in[`VWidth*(`APPRam_depth*23+7)-1:`VWidth*(`APPRam_depth*23+6)],data_in[`VWidth*(`APPRam_depth*22+7)-1:`VWidth*(`APPRam_depth*22+6)],data_in[`VWidth*(`APPRam_depth*21+7)-1:`VWidth*(`APPRam_depth*21+6)],data_in[`VWidth*(`APPRam_depth*20+7)-1:`VWidth*(`APPRam_depth*20+6)],data_in[`VWidth*(`APPRam_depth*19+7)-1:`VWidth*(`APPRam_depth*19+6)],data_in[`VWidth*(`APPRam_depth*18+7)-1:`VWidth*(`APPRam_depth*18+6)],data_in[`VWidth*(`APPRam_depth*17+7)-1:`VWidth*(`APPRam_depth*17+6)],data_in[`VWidth*(`APPRam_depth*16+7)-1:`VWidth*(`APPRam_depth*16+6)],data_in[`VWidth*(`APPRam_depth*15+7)-1:`VWidth*(`APPRam_depth*15+6)],data_in[`VWidth*(`APPRam_depth*14+7)-1:`VWidth*(`APPRam_depth*14+6)],data_in[`VWidth*(`APPRam_depth*13+7)-1:`VWidth*(`APPRam_depth*13+6)],data_in[`VWidth*(`APPRam_depth*12+7)-1:`VWidth*(`APPRam_depth*12+6)],data_in[`VWidth*(`APPRam_depth*11+7)-1:`VWidth*(`APPRam_depth*11+6)],data_in[`VWidth*(`APPRam_depth*10+7)-1:`VWidth*(`APPRam_depth*10+6)],data_in[`VWidth*(`APPRam_depth*9+7)-1:`VWidth*(`APPRam_depth*9+6)],data_in[`VWidth*(`APPRam_depth*8+7)-1:`VWidth*(`APPRam_depth*8+6)],data_in[`VWidth*(`APPRam_depth*7+7)-1:`VWidth*(`APPRam_depth*7+6)],data_in[`VWidth*(`APPRam_depth*6+7)-1:`VWidth*(`APPRam_depth*6+6)],data_in[`VWidth*(`APPRam_depth*5+7)-1:`VWidth*(`APPRam_depth*5+6)],data_in[`VWidth*(`APPRam_depth*4+7)-1:`VWidth*(`APPRam_depth*4+6)],data_in[`VWidth*(`APPRam_depth*3+7)-1:`VWidth*(`APPRam_depth*3+6)],data_in[`VWidth*(`APPRam_depth*2+7)-1:`VWidth*(`APPRam_depth*2+6)],data_in[`VWidth*(`APPRam_depth*1+7)-1:`VWidth*(`APPRam_depth*1+6)],data_in[`VWidth*(`APPRam_depth*0+7)-1:`VWidth*(`APPRam_depth*0+6)]};
			end
			7:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+8)-1:`VWidth*(`APPRam_depth*31+7)],data_in[`VWidth*(`APPRam_depth*30+8)-1:`VWidth*(`APPRam_depth*30+7)],data_in[`VWidth*(`APPRam_depth*29+8)-1:`VWidth*(`APPRam_depth*29+7)],data_in[`VWidth*(`APPRam_depth*28+8)-1:`VWidth*(`APPRam_depth*28+7)],data_in[`VWidth*(`APPRam_depth*27+8)-1:`VWidth*(`APPRam_depth*27+7)],data_in[`VWidth*(`APPRam_depth*26+8)-1:`VWidth*(`APPRam_depth*26+7)],data_in[`VWidth*(`APPRam_depth*25+8)-1:`VWidth*(`APPRam_depth*25+7)],data_in[`VWidth*(`APPRam_depth*24+8)-1:`VWidth*(`APPRam_depth*24+7)],data_in[`VWidth*(`APPRam_depth*23+8)-1:`VWidth*(`APPRam_depth*23+7)],data_in[`VWidth*(`APPRam_depth*22+8)-1:`VWidth*(`APPRam_depth*22+7)],data_in[`VWidth*(`APPRam_depth*21+8)-1:`VWidth*(`APPRam_depth*21+7)],data_in[`VWidth*(`APPRam_depth*20+8)-1:`VWidth*(`APPRam_depth*20+7)],data_in[`VWidth*(`APPRam_depth*19+8)-1:`VWidth*(`APPRam_depth*19+7)],data_in[`VWidth*(`APPRam_depth*18+8)-1:`VWidth*(`APPRam_depth*18+7)],data_in[`VWidth*(`APPRam_depth*17+8)-1:`VWidth*(`APPRam_depth*17+7)],data_in[`VWidth*(`APPRam_depth*16+8)-1:`VWidth*(`APPRam_depth*16+7)],data_in[`VWidth*(`APPRam_depth*15+8)-1:`VWidth*(`APPRam_depth*15+7)],data_in[`VWidth*(`APPRam_depth*14+8)-1:`VWidth*(`APPRam_depth*14+7)],data_in[`VWidth*(`APPRam_depth*13+8)-1:`VWidth*(`APPRam_depth*13+7)],data_in[`VWidth*(`APPRam_depth*12+8)-1:`VWidth*(`APPRam_depth*12+7)],data_in[`VWidth*(`APPRam_depth*11+8)-1:`VWidth*(`APPRam_depth*11+7)],data_in[`VWidth*(`APPRam_depth*10+8)-1:`VWidth*(`APPRam_depth*10+7)],data_in[`VWidth*(`APPRam_depth*9+8)-1:`VWidth*(`APPRam_depth*9+7)],data_in[`VWidth*(`APPRam_depth*8+8)-1:`VWidth*(`APPRam_depth*8+7)],data_in[`VWidth*(`APPRam_depth*7+8)-1:`VWidth*(`APPRam_depth*7+7)],data_in[`VWidth*(`APPRam_depth*6+8)-1:`VWidth*(`APPRam_depth*6+7)],data_in[`VWidth*(`APPRam_depth*5+8)-1:`VWidth*(`APPRam_depth*5+7)],data_in[`VWidth*(`APPRam_depth*4+8)-1:`VWidth*(`APPRam_depth*4+7)],data_in[`VWidth*(`APPRam_depth*3+8)-1:`VWidth*(`APPRam_depth*3+7)],data_in[`VWidth*(`APPRam_depth*2+8)-1:`VWidth*(`APPRam_depth*2+7)],data_in[`VWidth*(`APPRam_depth*1+8)-1:`VWidth*(`APPRam_depth*1+7)],data_in[`VWidth*(`APPRam_depth*0+8)-1:`VWidth*(`APPRam_depth*0+7)]};
			end
			8:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+9)-1:`VWidth*(`APPRam_depth*31+8)],data_in[`VWidth*(`APPRam_depth*30+9)-1:`VWidth*(`APPRam_depth*30+8)],data_in[`VWidth*(`APPRam_depth*29+9)-1:`VWidth*(`APPRam_depth*29+8)],data_in[`VWidth*(`APPRam_depth*28+9)-1:`VWidth*(`APPRam_depth*28+8)],data_in[`VWidth*(`APPRam_depth*27+9)-1:`VWidth*(`APPRam_depth*27+8)],data_in[`VWidth*(`APPRam_depth*26+9)-1:`VWidth*(`APPRam_depth*26+8)],data_in[`VWidth*(`APPRam_depth*25+9)-1:`VWidth*(`APPRam_depth*25+8)],data_in[`VWidth*(`APPRam_depth*24+9)-1:`VWidth*(`APPRam_depth*24+8)],data_in[`VWidth*(`APPRam_depth*23+9)-1:`VWidth*(`APPRam_depth*23+8)],data_in[`VWidth*(`APPRam_depth*22+9)-1:`VWidth*(`APPRam_depth*22+8)],data_in[`VWidth*(`APPRam_depth*21+9)-1:`VWidth*(`APPRam_depth*21+8)],data_in[`VWidth*(`APPRam_depth*20+9)-1:`VWidth*(`APPRam_depth*20+8)],data_in[`VWidth*(`APPRam_depth*19+9)-1:`VWidth*(`APPRam_depth*19+8)],data_in[`VWidth*(`APPRam_depth*18+9)-1:`VWidth*(`APPRam_depth*18+8)],data_in[`VWidth*(`APPRam_depth*17+9)-1:`VWidth*(`APPRam_depth*17+8)],data_in[`VWidth*(`APPRam_depth*16+9)-1:`VWidth*(`APPRam_depth*16+8)],data_in[`VWidth*(`APPRam_depth*15+9)-1:`VWidth*(`APPRam_depth*15+8)],data_in[`VWidth*(`APPRam_depth*14+9)-1:`VWidth*(`APPRam_depth*14+8)],data_in[`VWidth*(`APPRam_depth*13+9)-1:`VWidth*(`APPRam_depth*13+8)],data_in[`VWidth*(`APPRam_depth*12+9)-1:`VWidth*(`APPRam_depth*12+8)],data_in[`VWidth*(`APPRam_depth*11+9)-1:`VWidth*(`APPRam_depth*11+8)],data_in[`VWidth*(`APPRam_depth*10+9)-1:`VWidth*(`APPRam_depth*10+8)],data_in[`VWidth*(`APPRam_depth*9+9)-1:`VWidth*(`APPRam_depth*9+8)],data_in[`VWidth*(`APPRam_depth*8+9)-1:`VWidth*(`APPRam_depth*8+8)],data_in[`VWidth*(`APPRam_depth*7+9)-1:`VWidth*(`APPRam_depth*7+8)],data_in[`VWidth*(`APPRam_depth*6+9)-1:`VWidth*(`APPRam_depth*6+8)],data_in[`VWidth*(`APPRam_depth*5+9)-1:`VWidth*(`APPRam_depth*5+8)],data_in[`VWidth*(`APPRam_depth*4+9)-1:`VWidth*(`APPRam_depth*4+8)],data_in[`VWidth*(`APPRam_depth*3+9)-1:`VWidth*(`APPRam_depth*3+8)],data_in[`VWidth*(`APPRam_depth*2+9)-1:`VWidth*(`APPRam_depth*2+8)],data_in[`VWidth*(`APPRam_depth*1+9)-1:`VWidth*(`APPRam_depth*1+8)],data_in[`VWidth*(`APPRam_depth*0+9)-1:`VWidth*(`APPRam_depth*0+8)]};
			end
			9:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+10)-1:`VWidth*(`APPRam_depth*31+9)],data_in[`VWidth*(`APPRam_depth*30+10)-1:`VWidth*(`APPRam_depth*30+9)],data_in[`VWidth*(`APPRam_depth*29+10)-1:`VWidth*(`APPRam_depth*29+9)],data_in[`VWidth*(`APPRam_depth*28+10)-1:`VWidth*(`APPRam_depth*28+9)],data_in[`VWidth*(`APPRam_depth*27+10)-1:`VWidth*(`APPRam_depth*27+9)],data_in[`VWidth*(`APPRam_depth*26+10)-1:`VWidth*(`APPRam_depth*26+9)],data_in[`VWidth*(`APPRam_depth*25+10)-1:`VWidth*(`APPRam_depth*25+9)],data_in[`VWidth*(`APPRam_depth*24+10)-1:`VWidth*(`APPRam_depth*24+9)],data_in[`VWidth*(`APPRam_depth*23+10)-1:`VWidth*(`APPRam_depth*23+9)],data_in[`VWidth*(`APPRam_depth*22+10)-1:`VWidth*(`APPRam_depth*22+9)],data_in[`VWidth*(`APPRam_depth*21+10)-1:`VWidth*(`APPRam_depth*21+9)],data_in[`VWidth*(`APPRam_depth*20+10)-1:`VWidth*(`APPRam_depth*20+9)],data_in[`VWidth*(`APPRam_depth*19+10)-1:`VWidth*(`APPRam_depth*19+9)],data_in[`VWidth*(`APPRam_depth*18+10)-1:`VWidth*(`APPRam_depth*18+9)],data_in[`VWidth*(`APPRam_depth*17+10)-1:`VWidth*(`APPRam_depth*17+9)],data_in[`VWidth*(`APPRam_depth*16+10)-1:`VWidth*(`APPRam_depth*16+9)],data_in[`VWidth*(`APPRam_depth*15+10)-1:`VWidth*(`APPRam_depth*15+9)],data_in[`VWidth*(`APPRam_depth*14+10)-1:`VWidth*(`APPRam_depth*14+9)],data_in[`VWidth*(`APPRam_depth*13+10)-1:`VWidth*(`APPRam_depth*13+9)],data_in[`VWidth*(`APPRam_depth*12+10)-1:`VWidth*(`APPRam_depth*12+9)],data_in[`VWidth*(`APPRam_depth*11+10)-1:`VWidth*(`APPRam_depth*11+9)],data_in[`VWidth*(`APPRam_depth*10+10)-1:`VWidth*(`APPRam_depth*10+9)],data_in[`VWidth*(`APPRam_depth*9+10)-1:`VWidth*(`APPRam_depth*9+9)],data_in[`VWidth*(`APPRam_depth*8+10)-1:`VWidth*(`APPRam_depth*8+9)],data_in[`VWidth*(`APPRam_depth*7+10)-1:`VWidth*(`APPRam_depth*7+9)],data_in[`VWidth*(`APPRam_depth*6+10)-1:`VWidth*(`APPRam_depth*6+9)],data_in[`VWidth*(`APPRam_depth*5+10)-1:`VWidth*(`APPRam_depth*5+9)],data_in[`VWidth*(`APPRam_depth*4+10)-1:`VWidth*(`APPRam_depth*4+9)],data_in[`VWidth*(`APPRam_depth*3+10)-1:`VWidth*(`APPRam_depth*3+9)],data_in[`VWidth*(`APPRam_depth*2+10)-1:`VWidth*(`APPRam_depth*2+9)],data_in[`VWidth*(`APPRam_depth*1+10)-1:`VWidth*(`APPRam_depth*1+9)],data_in[`VWidth*(`APPRam_depth*0+10)-1:`VWidth*(`APPRam_depth*0+9)]};
			end
			10:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+11)-1:`VWidth*(`APPRam_depth*31+10)],data_in[`VWidth*(`APPRam_depth*30+11)-1:`VWidth*(`APPRam_depth*30+10)],data_in[`VWidth*(`APPRam_depth*29+11)-1:`VWidth*(`APPRam_depth*29+10)],data_in[`VWidth*(`APPRam_depth*28+11)-1:`VWidth*(`APPRam_depth*28+10)],data_in[`VWidth*(`APPRam_depth*27+11)-1:`VWidth*(`APPRam_depth*27+10)],data_in[`VWidth*(`APPRam_depth*26+11)-1:`VWidth*(`APPRam_depth*26+10)],data_in[`VWidth*(`APPRam_depth*25+11)-1:`VWidth*(`APPRam_depth*25+10)],data_in[`VWidth*(`APPRam_depth*24+11)-1:`VWidth*(`APPRam_depth*24+10)],data_in[`VWidth*(`APPRam_depth*23+11)-1:`VWidth*(`APPRam_depth*23+10)],data_in[`VWidth*(`APPRam_depth*22+11)-1:`VWidth*(`APPRam_depth*22+10)],data_in[`VWidth*(`APPRam_depth*21+11)-1:`VWidth*(`APPRam_depth*21+10)],data_in[`VWidth*(`APPRam_depth*20+11)-1:`VWidth*(`APPRam_depth*20+10)],data_in[`VWidth*(`APPRam_depth*19+11)-1:`VWidth*(`APPRam_depth*19+10)],data_in[`VWidth*(`APPRam_depth*18+11)-1:`VWidth*(`APPRam_depth*18+10)],data_in[`VWidth*(`APPRam_depth*17+11)-1:`VWidth*(`APPRam_depth*17+10)],data_in[`VWidth*(`APPRam_depth*16+11)-1:`VWidth*(`APPRam_depth*16+10)],data_in[`VWidth*(`APPRam_depth*15+11)-1:`VWidth*(`APPRam_depth*15+10)],data_in[`VWidth*(`APPRam_depth*14+11)-1:`VWidth*(`APPRam_depth*14+10)],data_in[`VWidth*(`APPRam_depth*13+11)-1:`VWidth*(`APPRam_depth*13+10)],data_in[`VWidth*(`APPRam_depth*12+11)-1:`VWidth*(`APPRam_depth*12+10)],data_in[`VWidth*(`APPRam_depth*11+11)-1:`VWidth*(`APPRam_depth*11+10)],data_in[`VWidth*(`APPRam_depth*10+11)-1:`VWidth*(`APPRam_depth*10+10)],data_in[`VWidth*(`APPRam_depth*9+11)-1:`VWidth*(`APPRam_depth*9+10)],data_in[`VWidth*(`APPRam_depth*8+11)-1:`VWidth*(`APPRam_depth*8+10)],data_in[`VWidth*(`APPRam_depth*7+11)-1:`VWidth*(`APPRam_depth*7+10)],data_in[`VWidth*(`APPRam_depth*6+11)-1:`VWidth*(`APPRam_depth*6+10)],data_in[`VWidth*(`APPRam_depth*5+11)-1:`VWidth*(`APPRam_depth*5+10)],data_in[`VWidth*(`APPRam_depth*4+11)-1:`VWidth*(`APPRam_depth*4+10)],data_in[`VWidth*(`APPRam_depth*3+11)-1:`VWidth*(`APPRam_depth*3+10)],data_in[`VWidth*(`APPRam_depth*2+11)-1:`VWidth*(`APPRam_depth*2+10)],data_in[`VWidth*(`APPRam_depth*1+11)-1:`VWidth*(`APPRam_depth*1+10)],data_in[`VWidth*(`APPRam_depth*0+11)-1:`VWidth*(`APPRam_depth*0+10)]};
			end
			11:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+12)-1:`VWidth*(`APPRam_depth*31+11)],data_in[`VWidth*(`APPRam_depth*30+12)-1:`VWidth*(`APPRam_depth*30+11)],data_in[`VWidth*(`APPRam_depth*29+12)-1:`VWidth*(`APPRam_depth*29+11)],data_in[`VWidth*(`APPRam_depth*28+12)-1:`VWidth*(`APPRam_depth*28+11)],data_in[`VWidth*(`APPRam_depth*27+12)-1:`VWidth*(`APPRam_depth*27+11)],data_in[`VWidth*(`APPRam_depth*26+12)-1:`VWidth*(`APPRam_depth*26+11)],data_in[`VWidth*(`APPRam_depth*25+12)-1:`VWidth*(`APPRam_depth*25+11)],data_in[`VWidth*(`APPRam_depth*24+12)-1:`VWidth*(`APPRam_depth*24+11)],data_in[`VWidth*(`APPRam_depth*23+12)-1:`VWidth*(`APPRam_depth*23+11)],data_in[`VWidth*(`APPRam_depth*22+12)-1:`VWidth*(`APPRam_depth*22+11)],data_in[`VWidth*(`APPRam_depth*21+12)-1:`VWidth*(`APPRam_depth*21+11)],data_in[`VWidth*(`APPRam_depth*20+12)-1:`VWidth*(`APPRam_depth*20+11)],data_in[`VWidth*(`APPRam_depth*19+12)-1:`VWidth*(`APPRam_depth*19+11)],data_in[`VWidth*(`APPRam_depth*18+12)-1:`VWidth*(`APPRam_depth*18+11)],data_in[`VWidth*(`APPRam_depth*17+12)-1:`VWidth*(`APPRam_depth*17+11)],data_in[`VWidth*(`APPRam_depth*16+12)-1:`VWidth*(`APPRam_depth*16+11)],data_in[`VWidth*(`APPRam_depth*15+12)-1:`VWidth*(`APPRam_depth*15+11)],data_in[`VWidth*(`APPRam_depth*14+12)-1:`VWidth*(`APPRam_depth*14+11)],data_in[`VWidth*(`APPRam_depth*13+12)-1:`VWidth*(`APPRam_depth*13+11)],data_in[`VWidth*(`APPRam_depth*12+12)-1:`VWidth*(`APPRam_depth*12+11)],data_in[`VWidth*(`APPRam_depth*11+12)-1:`VWidth*(`APPRam_depth*11+11)],data_in[`VWidth*(`APPRam_depth*10+12)-1:`VWidth*(`APPRam_depth*10+11)],data_in[`VWidth*(`APPRam_depth*9+12)-1:`VWidth*(`APPRam_depth*9+11)],data_in[`VWidth*(`APPRam_depth*8+12)-1:`VWidth*(`APPRam_depth*8+11)],data_in[`VWidth*(`APPRam_depth*7+12)-1:`VWidth*(`APPRam_depth*7+11)],data_in[`VWidth*(`APPRam_depth*6+12)-1:`VWidth*(`APPRam_depth*6+11)],data_in[`VWidth*(`APPRam_depth*5+12)-1:`VWidth*(`APPRam_depth*5+11)],data_in[`VWidth*(`APPRam_depth*4+12)-1:`VWidth*(`APPRam_depth*4+11)],data_in[`VWidth*(`APPRam_depth*3+12)-1:`VWidth*(`APPRam_depth*3+11)],data_in[`VWidth*(`APPRam_depth*2+12)-1:`VWidth*(`APPRam_depth*2+11)],data_in[`VWidth*(`APPRam_depth*1+12)-1:`VWidth*(`APPRam_depth*1+11)],data_in[`VWidth*(`APPRam_depth*0+12)-1:`VWidth*(`APPRam_depth*0+11)]};
			end
			12:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+13)-1:`VWidth*(`APPRam_depth*31+12)],data_in[`VWidth*(`APPRam_depth*30+13)-1:`VWidth*(`APPRam_depth*30+12)],data_in[`VWidth*(`APPRam_depth*29+13)-1:`VWidth*(`APPRam_depth*29+12)],data_in[`VWidth*(`APPRam_depth*28+13)-1:`VWidth*(`APPRam_depth*28+12)],data_in[`VWidth*(`APPRam_depth*27+13)-1:`VWidth*(`APPRam_depth*27+12)],data_in[`VWidth*(`APPRam_depth*26+13)-1:`VWidth*(`APPRam_depth*26+12)],data_in[`VWidth*(`APPRam_depth*25+13)-1:`VWidth*(`APPRam_depth*25+12)],data_in[`VWidth*(`APPRam_depth*24+13)-1:`VWidth*(`APPRam_depth*24+12)],data_in[`VWidth*(`APPRam_depth*23+13)-1:`VWidth*(`APPRam_depth*23+12)],data_in[`VWidth*(`APPRam_depth*22+13)-1:`VWidth*(`APPRam_depth*22+12)],data_in[`VWidth*(`APPRam_depth*21+13)-1:`VWidth*(`APPRam_depth*21+12)],data_in[`VWidth*(`APPRam_depth*20+13)-1:`VWidth*(`APPRam_depth*20+12)],data_in[`VWidth*(`APPRam_depth*19+13)-1:`VWidth*(`APPRam_depth*19+12)],data_in[`VWidth*(`APPRam_depth*18+13)-1:`VWidth*(`APPRam_depth*18+12)],data_in[`VWidth*(`APPRam_depth*17+13)-1:`VWidth*(`APPRam_depth*17+12)],data_in[`VWidth*(`APPRam_depth*16+13)-1:`VWidth*(`APPRam_depth*16+12)],data_in[`VWidth*(`APPRam_depth*15+13)-1:`VWidth*(`APPRam_depth*15+12)],data_in[`VWidth*(`APPRam_depth*14+13)-1:`VWidth*(`APPRam_depth*14+12)],data_in[`VWidth*(`APPRam_depth*13+13)-1:`VWidth*(`APPRam_depth*13+12)],data_in[`VWidth*(`APPRam_depth*12+13)-1:`VWidth*(`APPRam_depth*12+12)],data_in[`VWidth*(`APPRam_depth*11+13)-1:`VWidth*(`APPRam_depth*11+12)],data_in[`VWidth*(`APPRam_depth*10+13)-1:`VWidth*(`APPRam_depth*10+12)],data_in[`VWidth*(`APPRam_depth*9+13)-1:`VWidth*(`APPRam_depth*9+12)],data_in[`VWidth*(`APPRam_depth*8+13)-1:`VWidth*(`APPRam_depth*8+12)],data_in[`VWidth*(`APPRam_depth*7+13)-1:`VWidth*(`APPRam_depth*7+12)],data_in[`VWidth*(`APPRam_depth*6+13)-1:`VWidth*(`APPRam_depth*6+12)],data_in[`VWidth*(`APPRam_depth*5+13)-1:`VWidth*(`APPRam_depth*5+12)],data_in[`VWidth*(`APPRam_depth*4+13)-1:`VWidth*(`APPRam_depth*4+12)],data_in[`VWidth*(`APPRam_depth*3+13)-1:`VWidth*(`APPRam_depth*3+12)],data_in[`VWidth*(`APPRam_depth*2+13)-1:`VWidth*(`APPRam_depth*2+12)],data_in[`VWidth*(`APPRam_depth*1+13)-1:`VWidth*(`APPRam_depth*1+12)],data_in[`VWidth*(`APPRam_depth*0+13)-1:`VWidth*(`APPRam_depth*0+12)]};
			end
			13:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+14)-1:`VWidth*(`APPRam_depth*31+13)],data_in[`VWidth*(`APPRam_depth*30+14)-1:`VWidth*(`APPRam_depth*30+13)],data_in[`VWidth*(`APPRam_depth*29+14)-1:`VWidth*(`APPRam_depth*29+13)],data_in[`VWidth*(`APPRam_depth*28+14)-1:`VWidth*(`APPRam_depth*28+13)],data_in[`VWidth*(`APPRam_depth*27+14)-1:`VWidth*(`APPRam_depth*27+13)],data_in[`VWidth*(`APPRam_depth*26+14)-1:`VWidth*(`APPRam_depth*26+13)],data_in[`VWidth*(`APPRam_depth*25+14)-1:`VWidth*(`APPRam_depth*25+13)],data_in[`VWidth*(`APPRam_depth*24+14)-1:`VWidth*(`APPRam_depth*24+13)],data_in[`VWidth*(`APPRam_depth*23+14)-1:`VWidth*(`APPRam_depth*23+13)],data_in[`VWidth*(`APPRam_depth*22+14)-1:`VWidth*(`APPRam_depth*22+13)],data_in[`VWidth*(`APPRam_depth*21+14)-1:`VWidth*(`APPRam_depth*21+13)],data_in[`VWidth*(`APPRam_depth*20+14)-1:`VWidth*(`APPRam_depth*20+13)],data_in[`VWidth*(`APPRam_depth*19+14)-1:`VWidth*(`APPRam_depth*19+13)],data_in[`VWidth*(`APPRam_depth*18+14)-1:`VWidth*(`APPRam_depth*18+13)],data_in[`VWidth*(`APPRam_depth*17+14)-1:`VWidth*(`APPRam_depth*17+13)],data_in[`VWidth*(`APPRam_depth*16+14)-1:`VWidth*(`APPRam_depth*16+13)],data_in[`VWidth*(`APPRam_depth*15+14)-1:`VWidth*(`APPRam_depth*15+13)],data_in[`VWidth*(`APPRam_depth*14+14)-1:`VWidth*(`APPRam_depth*14+13)],data_in[`VWidth*(`APPRam_depth*13+14)-1:`VWidth*(`APPRam_depth*13+13)],data_in[`VWidth*(`APPRam_depth*12+14)-1:`VWidth*(`APPRam_depth*12+13)],data_in[`VWidth*(`APPRam_depth*11+14)-1:`VWidth*(`APPRam_depth*11+13)],data_in[`VWidth*(`APPRam_depth*10+14)-1:`VWidth*(`APPRam_depth*10+13)],data_in[`VWidth*(`APPRam_depth*9+14)-1:`VWidth*(`APPRam_depth*9+13)],data_in[`VWidth*(`APPRam_depth*8+14)-1:`VWidth*(`APPRam_depth*8+13)],data_in[`VWidth*(`APPRam_depth*7+14)-1:`VWidth*(`APPRam_depth*7+13)],data_in[`VWidth*(`APPRam_depth*6+14)-1:`VWidth*(`APPRam_depth*6+13)],data_in[`VWidth*(`APPRam_depth*5+14)-1:`VWidth*(`APPRam_depth*5+13)],data_in[`VWidth*(`APPRam_depth*4+14)-1:`VWidth*(`APPRam_depth*4+13)],data_in[`VWidth*(`APPRam_depth*3+14)-1:`VWidth*(`APPRam_depth*3+13)],data_in[`VWidth*(`APPRam_depth*2+14)-1:`VWidth*(`APPRam_depth*2+13)],data_in[`VWidth*(`APPRam_depth*1+14)-1:`VWidth*(`APPRam_depth*1+13)],data_in[`VWidth*(`APPRam_depth*0+14)-1:`VWidth*(`APPRam_depth*0+13)]};
			end
			14:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+15)-1:`VWidth*(`APPRam_depth*31+14)],data_in[`VWidth*(`APPRam_depth*30+15)-1:`VWidth*(`APPRam_depth*30+14)],data_in[`VWidth*(`APPRam_depth*29+15)-1:`VWidth*(`APPRam_depth*29+14)],data_in[`VWidth*(`APPRam_depth*28+15)-1:`VWidth*(`APPRam_depth*28+14)],data_in[`VWidth*(`APPRam_depth*27+15)-1:`VWidth*(`APPRam_depth*27+14)],data_in[`VWidth*(`APPRam_depth*26+15)-1:`VWidth*(`APPRam_depth*26+14)],data_in[`VWidth*(`APPRam_depth*25+15)-1:`VWidth*(`APPRam_depth*25+14)],data_in[`VWidth*(`APPRam_depth*24+15)-1:`VWidth*(`APPRam_depth*24+14)],data_in[`VWidth*(`APPRam_depth*23+15)-1:`VWidth*(`APPRam_depth*23+14)],data_in[`VWidth*(`APPRam_depth*22+15)-1:`VWidth*(`APPRam_depth*22+14)],data_in[`VWidth*(`APPRam_depth*21+15)-1:`VWidth*(`APPRam_depth*21+14)],data_in[`VWidth*(`APPRam_depth*20+15)-1:`VWidth*(`APPRam_depth*20+14)],data_in[`VWidth*(`APPRam_depth*19+15)-1:`VWidth*(`APPRam_depth*19+14)],data_in[`VWidth*(`APPRam_depth*18+15)-1:`VWidth*(`APPRam_depth*18+14)],data_in[`VWidth*(`APPRam_depth*17+15)-1:`VWidth*(`APPRam_depth*17+14)],data_in[`VWidth*(`APPRam_depth*16+15)-1:`VWidth*(`APPRam_depth*16+14)],data_in[`VWidth*(`APPRam_depth*15+15)-1:`VWidth*(`APPRam_depth*15+14)],data_in[`VWidth*(`APPRam_depth*14+15)-1:`VWidth*(`APPRam_depth*14+14)],data_in[`VWidth*(`APPRam_depth*13+15)-1:`VWidth*(`APPRam_depth*13+14)],data_in[`VWidth*(`APPRam_depth*12+15)-1:`VWidth*(`APPRam_depth*12+14)],data_in[`VWidth*(`APPRam_depth*11+15)-1:`VWidth*(`APPRam_depth*11+14)],data_in[`VWidth*(`APPRam_depth*10+15)-1:`VWidth*(`APPRam_depth*10+14)],data_in[`VWidth*(`APPRam_depth*9+15)-1:`VWidth*(`APPRam_depth*9+14)],data_in[`VWidth*(`APPRam_depth*8+15)-1:`VWidth*(`APPRam_depth*8+14)],data_in[`VWidth*(`APPRam_depth*7+15)-1:`VWidth*(`APPRam_depth*7+14)],data_in[`VWidth*(`APPRam_depth*6+15)-1:`VWidth*(`APPRam_depth*6+14)],data_in[`VWidth*(`APPRam_depth*5+15)-1:`VWidth*(`APPRam_depth*5+14)],data_in[`VWidth*(`APPRam_depth*4+15)-1:`VWidth*(`APPRam_depth*4+14)],data_in[`VWidth*(`APPRam_depth*3+15)-1:`VWidth*(`APPRam_depth*3+14)],data_in[`VWidth*(`APPRam_depth*2+15)-1:`VWidth*(`APPRam_depth*2+14)],data_in[`VWidth*(`APPRam_depth*1+15)-1:`VWidth*(`APPRam_depth*1+14)],data_in[`VWidth*(`APPRam_depth*0+15)-1:`VWidth*(`APPRam_depth*0+14)]};
			end
			15:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+16)-1:`VWidth*(`APPRam_depth*31+15)],data_in[`VWidth*(`APPRam_depth*30+16)-1:`VWidth*(`APPRam_depth*30+15)],data_in[`VWidth*(`APPRam_depth*29+16)-1:`VWidth*(`APPRam_depth*29+15)],data_in[`VWidth*(`APPRam_depth*28+16)-1:`VWidth*(`APPRam_depth*28+15)],data_in[`VWidth*(`APPRam_depth*27+16)-1:`VWidth*(`APPRam_depth*27+15)],data_in[`VWidth*(`APPRam_depth*26+16)-1:`VWidth*(`APPRam_depth*26+15)],data_in[`VWidth*(`APPRam_depth*25+16)-1:`VWidth*(`APPRam_depth*25+15)],data_in[`VWidth*(`APPRam_depth*24+16)-1:`VWidth*(`APPRam_depth*24+15)],data_in[`VWidth*(`APPRam_depth*23+16)-1:`VWidth*(`APPRam_depth*23+15)],data_in[`VWidth*(`APPRam_depth*22+16)-1:`VWidth*(`APPRam_depth*22+15)],data_in[`VWidth*(`APPRam_depth*21+16)-1:`VWidth*(`APPRam_depth*21+15)],data_in[`VWidth*(`APPRam_depth*20+16)-1:`VWidth*(`APPRam_depth*20+15)],data_in[`VWidth*(`APPRam_depth*19+16)-1:`VWidth*(`APPRam_depth*19+15)],data_in[`VWidth*(`APPRam_depth*18+16)-1:`VWidth*(`APPRam_depth*18+15)],data_in[`VWidth*(`APPRam_depth*17+16)-1:`VWidth*(`APPRam_depth*17+15)],data_in[`VWidth*(`APPRam_depth*16+16)-1:`VWidth*(`APPRam_depth*16+15)],data_in[`VWidth*(`APPRam_depth*15+16)-1:`VWidth*(`APPRam_depth*15+15)],data_in[`VWidth*(`APPRam_depth*14+16)-1:`VWidth*(`APPRam_depth*14+15)],data_in[`VWidth*(`APPRam_depth*13+16)-1:`VWidth*(`APPRam_depth*13+15)],data_in[`VWidth*(`APPRam_depth*12+16)-1:`VWidth*(`APPRam_depth*12+15)],data_in[`VWidth*(`APPRam_depth*11+16)-1:`VWidth*(`APPRam_depth*11+15)],data_in[`VWidth*(`APPRam_depth*10+16)-1:`VWidth*(`APPRam_depth*10+15)],data_in[`VWidth*(`APPRam_depth*9+16)-1:`VWidth*(`APPRam_depth*9+15)],data_in[`VWidth*(`APPRam_depth*8+16)-1:`VWidth*(`APPRam_depth*8+15)],data_in[`VWidth*(`APPRam_depth*7+16)-1:`VWidth*(`APPRam_depth*7+15)],data_in[`VWidth*(`APPRam_depth*6+16)-1:`VWidth*(`APPRam_depth*6+15)],data_in[`VWidth*(`APPRam_depth*5+16)-1:`VWidth*(`APPRam_depth*5+15)],data_in[`VWidth*(`APPRam_depth*4+16)-1:`VWidth*(`APPRam_depth*4+15)],data_in[`VWidth*(`APPRam_depth*3+16)-1:`VWidth*(`APPRam_depth*3+15)],data_in[`VWidth*(`APPRam_depth*2+16)-1:`VWidth*(`APPRam_depth*2+15)],data_in[`VWidth*(`APPRam_depth*1+16)-1:`VWidth*(`APPRam_depth*1+15)],data_in[`VWidth*(`APPRam_depth*0+16)-1:`VWidth*(`APPRam_depth*0+15)]};
			end
			16:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+17)-1:`VWidth*(`APPRam_depth*31+16)],data_in[`VWidth*(`APPRam_depth*30+17)-1:`VWidth*(`APPRam_depth*30+16)],data_in[`VWidth*(`APPRam_depth*29+17)-1:`VWidth*(`APPRam_depth*29+16)],data_in[`VWidth*(`APPRam_depth*28+17)-1:`VWidth*(`APPRam_depth*28+16)],data_in[`VWidth*(`APPRam_depth*27+17)-1:`VWidth*(`APPRam_depth*27+16)],data_in[`VWidth*(`APPRam_depth*26+17)-1:`VWidth*(`APPRam_depth*26+16)],data_in[`VWidth*(`APPRam_depth*25+17)-1:`VWidth*(`APPRam_depth*25+16)],data_in[`VWidth*(`APPRam_depth*24+17)-1:`VWidth*(`APPRam_depth*24+16)],data_in[`VWidth*(`APPRam_depth*23+17)-1:`VWidth*(`APPRam_depth*23+16)],data_in[`VWidth*(`APPRam_depth*22+17)-1:`VWidth*(`APPRam_depth*22+16)],data_in[`VWidth*(`APPRam_depth*21+17)-1:`VWidth*(`APPRam_depth*21+16)],data_in[`VWidth*(`APPRam_depth*20+17)-1:`VWidth*(`APPRam_depth*20+16)],data_in[`VWidth*(`APPRam_depth*19+17)-1:`VWidth*(`APPRam_depth*19+16)],data_in[`VWidth*(`APPRam_depth*18+17)-1:`VWidth*(`APPRam_depth*18+16)],data_in[`VWidth*(`APPRam_depth*17+17)-1:`VWidth*(`APPRam_depth*17+16)],data_in[`VWidth*(`APPRam_depth*16+17)-1:`VWidth*(`APPRam_depth*16+16)],data_in[`VWidth*(`APPRam_depth*15+17)-1:`VWidth*(`APPRam_depth*15+16)],data_in[`VWidth*(`APPRam_depth*14+17)-1:`VWidth*(`APPRam_depth*14+16)],data_in[`VWidth*(`APPRam_depth*13+17)-1:`VWidth*(`APPRam_depth*13+16)],data_in[`VWidth*(`APPRam_depth*12+17)-1:`VWidth*(`APPRam_depth*12+16)],data_in[`VWidth*(`APPRam_depth*11+17)-1:`VWidth*(`APPRam_depth*11+16)],data_in[`VWidth*(`APPRam_depth*10+17)-1:`VWidth*(`APPRam_depth*10+16)],data_in[`VWidth*(`APPRam_depth*9+17)-1:`VWidth*(`APPRam_depth*9+16)],data_in[`VWidth*(`APPRam_depth*8+17)-1:`VWidth*(`APPRam_depth*8+16)],data_in[`VWidth*(`APPRam_depth*7+17)-1:`VWidth*(`APPRam_depth*7+16)],data_in[`VWidth*(`APPRam_depth*6+17)-1:`VWidth*(`APPRam_depth*6+16)],data_in[`VWidth*(`APPRam_depth*5+17)-1:`VWidth*(`APPRam_depth*5+16)],data_in[`VWidth*(`APPRam_depth*4+17)-1:`VWidth*(`APPRam_depth*4+16)],data_in[`VWidth*(`APPRam_depth*3+17)-1:`VWidth*(`APPRam_depth*3+16)],data_in[`VWidth*(`APPRam_depth*2+17)-1:`VWidth*(`APPRam_depth*2+16)],data_in[`VWidth*(`APPRam_depth*1+17)-1:`VWidth*(`APPRam_depth*1+16)],data_in[`VWidth*(`APPRam_depth*0+17)-1:`VWidth*(`APPRam_depth*0+16)]};
			end
			17:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+18)-1:`VWidth*(`APPRam_depth*31+17)],data_in[`VWidth*(`APPRam_depth*30+18)-1:`VWidth*(`APPRam_depth*30+17)],data_in[`VWidth*(`APPRam_depth*29+18)-1:`VWidth*(`APPRam_depth*29+17)],data_in[`VWidth*(`APPRam_depth*28+18)-1:`VWidth*(`APPRam_depth*28+17)],data_in[`VWidth*(`APPRam_depth*27+18)-1:`VWidth*(`APPRam_depth*27+17)],data_in[`VWidth*(`APPRam_depth*26+18)-1:`VWidth*(`APPRam_depth*26+17)],data_in[`VWidth*(`APPRam_depth*25+18)-1:`VWidth*(`APPRam_depth*25+17)],data_in[`VWidth*(`APPRam_depth*24+18)-1:`VWidth*(`APPRam_depth*24+17)],data_in[`VWidth*(`APPRam_depth*23+18)-1:`VWidth*(`APPRam_depth*23+17)],data_in[`VWidth*(`APPRam_depth*22+18)-1:`VWidth*(`APPRam_depth*22+17)],data_in[`VWidth*(`APPRam_depth*21+18)-1:`VWidth*(`APPRam_depth*21+17)],data_in[`VWidth*(`APPRam_depth*20+18)-1:`VWidth*(`APPRam_depth*20+17)],data_in[`VWidth*(`APPRam_depth*19+18)-1:`VWidth*(`APPRam_depth*19+17)],data_in[`VWidth*(`APPRam_depth*18+18)-1:`VWidth*(`APPRam_depth*18+17)],data_in[`VWidth*(`APPRam_depth*17+18)-1:`VWidth*(`APPRam_depth*17+17)],data_in[`VWidth*(`APPRam_depth*16+18)-1:`VWidth*(`APPRam_depth*16+17)],data_in[`VWidth*(`APPRam_depth*15+18)-1:`VWidth*(`APPRam_depth*15+17)],data_in[`VWidth*(`APPRam_depth*14+18)-1:`VWidth*(`APPRam_depth*14+17)],data_in[`VWidth*(`APPRam_depth*13+18)-1:`VWidth*(`APPRam_depth*13+17)],data_in[`VWidth*(`APPRam_depth*12+18)-1:`VWidth*(`APPRam_depth*12+17)],data_in[`VWidth*(`APPRam_depth*11+18)-1:`VWidth*(`APPRam_depth*11+17)],data_in[`VWidth*(`APPRam_depth*10+18)-1:`VWidth*(`APPRam_depth*10+17)],data_in[`VWidth*(`APPRam_depth*9+18)-1:`VWidth*(`APPRam_depth*9+17)],data_in[`VWidth*(`APPRam_depth*8+18)-1:`VWidth*(`APPRam_depth*8+17)],data_in[`VWidth*(`APPRam_depth*7+18)-1:`VWidth*(`APPRam_depth*7+17)],data_in[`VWidth*(`APPRam_depth*6+18)-1:`VWidth*(`APPRam_depth*6+17)],data_in[`VWidth*(`APPRam_depth*5+18)-1:`VWidth*(`APPRam_depth*5+17)],data_in[`VWidth*(`APPRam_depth*4+18)-1:`VWidth*(`APPRam_depth*4+17)],data_in[`VWidth*(`APPRam_depth*3+18)-1:`VWidth*(`APPRam_depth*3+17)],data_in[`VWidth*(`APPRam_depth*2+18)-1:`VWidth*(`APPRam_depth*2+17)],data_in[`VWidth*(`APPRam_depth*1+18)-1:`VWidth*(`APPRam_depth*1+17)],data_in[`VWidth*(`APPRam_depth*0+18)-1:`VWidth*(`APPRam_depth*0+17)]};
			end
			18:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+19)-1:`VWidth*(`APPRam_depth*31+18)],data_in[`VWidth*(`APPRam_depth*30+19)-1:`VWidth*(`APPRam_depth*30+18)],data_in[`VWidth*(`APPRam_depth*29+19)-1:`VWidth*(`APPRam_depth*29+18)],data_in[`VWidth*(`APPRam_depth*28+19)-1:`VWidth*(`APPRam_depth*28+18)],data_in[`VWidth*(`APPRam_depth*27+19)-1:`VWidth*(`APPRam_depth*27+18)],data_in[`VWidth*(`APPRam_depth*26+19)-1:`VWidth*(`APPRam_depth*26+18)],data_in[`VWidth*(`APPRam_depth*25+19)-1:`VWidth*(`APPRam_depth*25+18)],data_in[`VWidth*(`APPRam_depth*24+19)-1:`VWidth*(`APPRam_depth*24+18)],data_in[`VWidth*(`APPRam_depth*23+19)-1:`VWidth*(`APPRam_depth*23+18)],data_in[`VWidth*(`APPRam_depth*22+19)-1:`VWidth*(`APPRam_depth*22+18)],data_in[`VWidth*(`APPRam_depth*21+19)-1:`VWidth*(`APPRam_depth*21+18)],data_in[`VWidth*(`APPRam_depth*20+19)-1:`VWidth*(`APPRam_depth*20+18)],data_in[`VWidth*(`APPRam_depth*19+19)-1:`VWidth*(`APPRam_depth*19+18)],data_in[`VWidth*(`APPRam_depth*18+19)-1:`VWidth*(`APPRam_depth*18+18)],data_in[`VWidth*(`APPRam_depth*17+19)-1:`VWidth*(`APPRam_depth*17+18)],data_in[`VWidth*(`APPRam_depth*16+19)-1:`VWidth*(`APPRam_depth*16+18)],data_in[`VWidth*(`APPRam_depth*15+19)-1:`VWidth*(`APPRam_depth*15+18)],data_in[`VWidth*(`APPRam_depth*14+19)-1:`VWidth*(`APPRam_depth*14+18)],data_in[`VWidth*(`APPRam_depth*13+19)-1:`VWidth*(`APPRam_depth*13+18)],data_in[`VWidth*(`APPRam_depth*12+19)-1:`VWidth*(`APPRam_depth*12+18)],data_in[`VWidth*(`APPRam_depth*11+19)-1:`VWidth*(`APPRam_depth*11+18)],data_in[`VWidth*(`APPRam_depth*10+19)-1:`VWidth*(`APPRam_depth*10+18)],data_in[`VWidth*(`APPRam_depth*9+19)-1:`VWidth*(`APPRam_depth*9+18)],data_in[`VWidth*(`APPRam_depth*8+19)-1:`VWidth*(`APPRam_depth*8+18)],data_in[`VWidth*(`APPRam_depth*7+19)-1:`VWidth*(`APPRam_depth*7+18)],data_in[`VWidth*(`APPRam_depth*6+19)-1:`VWidth*(`APPRam_depth*6+18)],data_in[`VWidth*(`APPRam_depth*5+19)-1:`VWidth*(`APPRam_depth*5+18)],data_in[`VWidth*(`APPRam_depth*4+19)-1:`VWidth*(`APPRam_depth*4+18)],data_in[`VWidth*(`APPRam_depth*3+19)-1:`VWidth*(`APPRam_depth*3+18)],data_in[`VWidth*(`APPRam_depth*2+19)-1:`VWidth*(`APPRam_depth*2+18)],data_in[`VWidth*(`APPRam_depth*1+19)-1:`VWidth*(`APPRam_depth*1+18)],data_in[`VWidth*(`APPRam_depth*0+19)-1:`VWidth*(`APPRam_depth*0+18)]};
			end
			19:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+20)-1:`VWidth*(`APPRam_depth*31+19)],data_in[`VWidth*(`APPRam_depth*30+20)-1:`VWidth*(`APPRam_depth*30+19)],data_in[`VWidth*(`APPRam_depth*29+20)-1:`VWidth*(`APPRam_depth*29+19)],data_in[`VWidth*(`APPRam_depth*28+20)-1:`VWidth*(`APPRam_depth*28+19)],data_in[`VWidth*(`APPRam_depth*27+20)-1:`VWidth*(`APPRam_depth*27+19)],data_in[`VWidth*(`APPRam_depth*26+20)-1:`VWidth*(`APPRam_depth*26+19)],data_in[`VWidth*(`APPRam_depth*25+20)-1:`VWidth*(`APPRam_depth*25+19)],data_in[`VWidth*(`APPRam_depth*24+20)-1:`VWidth*(`APPRam_depth*24+19)],data_in[`VWidth*(`APPRam_depth*23+20)-1:`VWidth*(`APPRam_depth*23+19)],data_in[`VWidth*(`APPRam_depth*22+20)-1:`VWidth*(`APPRam_depth*22+19)],data_in[`VWidth*(`APPRam_depth*21+20)-1:`VWidth*(`APPRam_depth*21+19)],data_in[`VWidth*(`APPRam_depth*20+20)-1:`VWidth*(`APPRam_depth*20+19)],data_in[`VWidth*(`APPRam_depth*19+20)-1:`VWidth*(`APPRam_depth*19+19)],data_in[`VWidth*(`APPRam_depth*18+20)-1:`VWidth*(`APPRam_depth*18+19)],data_in[`VWidth*(`APPRam_depth*17+20)-1:`VWidth*(`APPRam_depth*17+19)],data_in[`VWidth*(`APPRam_depth*16+20)-1:`VWidth*(`APPRam_depth*16+19)],data_in[`VWidth*(`APPRam_depth*15+20)-1:`VWidth*(`APPRam_depth*15+19)],data_in[`VWidth*(`APPRam_depth*14+20)-1:`VWidth*(`APPRam_depth*14+19)],data_in[`VWidth*(`APPRam_depth*13+20)-1:`VWidth*(`APPRam_depth*13+19)],data_in[`VWidth*(`APPRam_depth*12+20)-1:`VWidth*(`APPRam_depth*12+19)],data_in[`VWidth*(`APPRam_depth*11+20)-1:`VWidth*(`APPRam_depth*11+19)],data_in[`VWidth*(`APPRam_depth*10+20)-1:`VWidth*(`APPRam_depth*10+19)],data_in[`VWidth*(`APPRam_depth*9+20)-1:`VWidth*(`APPRam_depth*9+19)],data_in[`VWidth*(`APPRam_depth*8+20)-1:`VWidth*(`APPRam_depth*8+19)],data_in[`VWidth*(`APPRam_depth*7+20)-1:`VWidth*(`APPRam_depth*7+19)],data_in[`VWidth*(`APPRam_depth*6+20)-1:`VWidth*(`APPRam_depth*6+19)],data_in[`VWidth*(`APPRam_depth*5+20)-1:`VWidth*(`APPRam_depth*5+19)],data_in[`VWidth*(`APPRam_depth*4+20)-1:`VWidth*(`APPRam_depth*4+19)],data_in[`VWidth*(`APPRam_depth*3+20)-1:`VWidth*(`APPRam_depth*3+19)],data_in[`VWidth*(`APPRam_depth*2+20)-1:`VWidth*(`APPRam_depth*2+19)],data_in[`VWidth*(`APPRam_depth*1+20)-1:`VWidth*(`APPRam_depth*1+19)],data_in[`VWidth*(`APPRam_depth*0+20)-1:`VWidth*(`APPRam_depth*0+19)]};
			end
			20:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+21)-1:`VWidth*(`APPRam_depth*31+20)],data_in[`VWidth*(`APPRam_depth*30+21)-1:`VWidth*(`APPRam_depth*30+20)],data_in[`VWidth*(`APPRam_depth*29+21)-1:`VWidth*(`APPRam_depth*29+20)],data_in[`VWidth*(`APPRam_depth*28+21)-1:`VWidth*(`APPRam_depth*28+20)],data_in[`VWidth*(`APPRam_depth*27+21)-1:`VWidth*(`APPRam_depth*27+20)],data_in[`VWidth*(`APPRam_depth*26+21)-1:`VWidth*(`APPRam_depth*26+20)],data_in[`VWidth*(`APPRam_depth*25+21)-1:`VWidth*(`APPRam_depth*25+20)],data_in[`VWidth*(`APPRam_depth*24+21)-1:`VWidth*(`APPRam_depth*24+20)],data_in[`VWidth*(`APPRam_depth*23+21)-1:`VWidth*(`APPRam_depth*23+20)],data_in[`VWidth*(`APPRam_depth*22+21)-1:`VWidth*(`APPRam_depth*22+20)],data_in[`VWidth*(`APPRam_depth*21+21)-1:`VWidth*(`APPRam_depth*21+20)],data_in[`VWidth*(`APPRam_depth*20+21)-1:`VWidth*(`APPRam_depth*20+20)],data_in[`VWidth*(`APPRam_depth*19+21)-1:`VWidth*(`APPRam_depth*19+20)],data_in[`VWidth*(`APPRam_depth*18+21)-1:`VWidth*(`APPRam_depth*18+20)],data_in[`VWidth*(`APPRam_depth*17+21)-1:`VWidth*(`APPRam_depth*17+20)],data_in[`VWidth*(`APPRam_depth*16+21)-1:`VWidth*(`APPRam_depth*16+20)],data_in[`VWidth*(`APPRam_depth*15+21)-1:`VWidth*(`APPRam_depth*15+20)],data_in[`VWidth*(`APPRam_depth*14+21)-1:`VWidth*(`APPRam_depth*14+20)],data_in[`VWidth*(`APPRam_depth*13+21)-1:`VWidth*(`APPRam_depth*13+20)],data_in[`VWidth*(`APPRam_depth*12+21)-1:`VWidth*(`APPRam_depth*12+20)],data_in[`VWidth*(`APPRam_depth*11+21)-1:`VWidth*(`APPRam_depth*11+20)],data_in[`VWidth*(`APPRam_depth*10+21)-1:`VWidth*(`APPRam_depth*10+20)],data_in[`VWidth*(`APPRam_depth*9+21)-1:`VWidth*(`APPRam_depth*9+20)],data_in[`VWidth*(`APPRam_depth*8+21)-1:`VWidth*(`APPRam_depth*8+20)],data_in[`VWidth*(`APPRam_depth*7+21)-1:`VWidth*(`APPRam_depth*7+20)],data_in[`VWidth*(`APPRam_depth*6+21)-1:`VWidth*(`APPRam_depth*6+20)],data_in[`VWidth*(`APPRam_depth*5+21)-1:`VWidth*(`APPRam_depth*5+20)],data_in[`VWidth*(`APPRam_depth*4+21)-1:`VWidth*(`APPRam_depth*4+20)],data_in[`VWidth*(`APPRam_depth*3+21)-1:`VWidth*(`APPRam_depth*3+20)],data_in[`VWidth*(`APPRam_depth*2+21)-1:`VWidth*(`APPRam_depth*2+20)],data_in[`VWidth*(`APPRam_depth*1+21)-1:`VWidth*(`APPRam_depth*1+20)],data_in[`VWidth*(`APPRam_depth*0+21)-1:`VWidth*(`APPRam_depth*0+20)]};
			end
			21:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+22)-1:`VWidth*(`APPRam_depth*31+21)],data_in[`VWidth*(`APPRam_depth*30+22)-1:`VWidth*(`APPRam_depth*30+21)],data_in[`VWidth*(`APPRam_depth*29+22)-1:`VWidth*(`APPRam_depth*29+21)],data_in[`VWidth*(`APPRam_depth*28+22)-1:`VWidth*(`APPRam_depth*28+21)],data_in[`VWidth*(`APPRam_depth*27+22)-1:`VWidth*(`APPRam_depth*27+21)],data_in[`VWidth*(`APPRam_depth*26+22)-1:`VWidth*(`APPRam_depth*26+21)],data_in[`VWidth*(`APPRam_depth*25+22)-1:`VWidth*(`APPRam_depth*25+21)],data_in[`VWidth*(`APPRam_depth*24+22)-1:`VWidth*(`APPRam_depth*24+21)],data_in[`VWidth*(`APPRam_depth*23+22)-1:`VWidth*(`APPRam_depth*23+21)],data_in[`VWidth*(`APPRam_depth*22+22)-1:`VWidth*(`APPRam_depth*22+21)],data_in[`VWidth*(`APPRam_depth*21+22)-1:`VWidth*(`APPRam_depth*21+21)],data_in[`VWidth*(`APPRam_depth*20+22)-1:`VWidth*(`APPRam_depth*20+21)],data_in[`VWidth*(`APPRam_depth*19+22)-1:`VWidth*(`APPRam_depth*19+21)],data_in[`VWidth*(`APPRam_depth*18+22)-1:`VWidth*(`APPRam_depth*18+21)],data_in[`VWidth*(`APPRam_depth*17+22)-1:`VWidth*(`APPRam_depth*17+21)],data_in[`VWidth*(`APPRam_depth*16+22)-1:`VWidth*(`APPRam_depth*16+21)],data_in[`VWidth*(`APPRam_depth*15+22)-1:`VWidth*(`APPRam_depth*15+21)],data_in[`VWidth*(`APPRam_depth*14+22)-1:`VWidth*(`APPRam_depth*14+21)],data_in[`VWidth*(`APPRam_depth*13+22)-1:`VWidth*(`APPRam_depth*13+21)],data_in[`VWidth*(`APPRam_depth*12+22)-1:`VWidth*(`APPRam_depth*12+21)],data_in[`VWidth*(`APPRam_depth*11+22)-1:`VWidth*(`APPRam_depth*11+21)],data_in[`VWidth*(`APPRam_depth*10+22)-1:`VWidth*(`APPRam_depth*10+21)],data_in[`VWidth*(`APPRam_depth*9+22)-1:`VWidth*(`APPRam_depth*9+21)],data_in[`VWidth*(`APPRam_depth*8+22)-1:`VWidth*(`APPRam_depth*8+21)],data_in[`VWidth*(`APPRam_depth*7+22)-1:`VWidth*(`APPRam_depth*7+21)],data_in[`VWidth*(`APPRam_depth*6+22)-1:`VWidth*(`APPRam_depth*6+21)],data_in[`VWidth*(`APPRam_depth*5+22)-1:`VWidth*(`APPRam_depth*5+21)],data_in[`VWidth*(`APPRam_depth*4+22)-1:`VWidth*(`APPRam_depth*4+21)],data_in[`VWidth*(`APPRam_depth*3+22)-1:`VWidth*(`APPRam_depth*3+21)],data_in[`VWidth*(`APPRam_depth*2+22)-1:`VWidth*(`APPRam_depth*2+21)],data_in[`VWidth*(`APPRam_depth*1+22)-1:`VWidth*(`APPRam_depth*1+21)],data_in[`VWidth*(`APPRam_depth*0+22)-1:`VWidth*(`APPRam_depth*0+21)]};
			end
			22:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+23)-1:`VWidth*(`APPRam_depth*31+22)],data_in[`VWidth*(`APPRam_depth*30+23)-1:`VWidth*(`APPRam_depth*30+22)],data_in[`VWidth*(`APPRam_depth*29+23)-1:`VWidth*(`APPRam_depth*29+22)],data_in[`VWidth*(`APPRam_depth*28+23)-1:`VWidth*(`APPRam_depth*28+22)],data_in[`VWidth*(`APPRam_depth*27+23)-1:`VWidth*(`APPRam_depth*27+22)],data_in[`VWidth*(`APPRam_depth*26+23)-1:`VWidth*(`APPRam_depth*26+22)],data_in[`VWidth*(`APPRam_depth*25+23)-1:`VWidth*(`APPRam_depth*25+22)],data_in[`VWidth*(`APPRam_depth*24+23)-1:`VWidth*(`APPRam_depth*24+22)],data_in[`VWidth*(`APPRam_depth*23+23)-1:`VWidth*(`APPRam_depth*23+22)],data_in[`VWidth*(`APPRam_depth*22+23)-1:`VWidth*(`APPRam_depth*22+22)],data_in[`VWidth*(`APPRam_depth*21+23)-1:`VWidth*(`APPRam_depth*21+22)],data_in[`VWidth*(`APPRam_depth*20+23)-1:`VWidth*(`APPRam_depth*20+22)],data_in[`VWidth*(`APPRam_depth*19+23)-1:`VWidth*(`APPRam_depth*19+22)],data_in[`VWidth*(`APPRam_depth*18+23)-1:`VWidth*(`APPRam_depth*18+22)],data_in[`VWidth*(`APPRam_depth*17+23)-1:`VWidth*(`APPRam_depth*17+22)],data_in[`VWidth*(`APPRam_depth*16+23)-1:`VWidth*(`APPRam_depth*16+22)],data_in[`VWidth*(`APPRam_depth*15+23)-1:`VWidth*(`APPRam_depth*15+22)],data_in[`VWidth*(`APPRam_depth*14+23)-1:`VWidth*(`APPRam_depth*14+22)],data_in[`VWidth*(`APPRam_depth*13+23)-1:`VWidth*(`APPRam_depth*13+22)],data_in[`VWidth*(`APPRam_depth*12+23)-1:`VWidth*(`APPRam_depth*12+22)],data_in[`VWidth*(`APPRam_depth*11+23)-1:`VWidth*(`APPRam_depth*11+22)],data_in[`VWidth*(`APPRam_depth*10+23)-1:`VWidth*(`APPRam_depth*10+22)],data_in[`VWidth*(`APPRam_depth*9+23)-1:`VWidth*(`APPRam_depth*9+22)],data_in[`VWidth*(`APPRam_depth*8+23)-1:`VWidth*(`APPRam_depth*8+22)],data_in[`VWidth*(`APPRam_depth*7+23)-1:`VWidth*(`APPRam_depth*7+22)],data_in[`VWidth*(`APPRam_depth*6+23)-1:`VWidth*(`APPRam_depth*6+22)],data_in[`VWidth*(`APPRam_depth*5+23)-1:`VWidth*(`APPRam_depth*5+22)],data_in[`VWidth*(`APPRam_depth*4+23)-1:`VWidth*(`APPRam_depth*4+22)],data_in[`VWidth*(`APPRam_depth*3+23)-1:`VWidth*(`APPRam_depth*3+22)],data_in[`VWidth*(`APPRam_depth*2+23)-1:`VWidth*(`APPRam_depth*2+22)],data_in[`VWidth*(`APPRam_depth*1+23)-1:`VWidth*(`APPRam_depth*1+22)],data_in[`VWidth*(`APPRam_depth*0+23)-1:`VWidth*(`APPRam_depth*0+22)]};
			end
			23:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+24)-1:`VWidth*(`APPRam_depth*31+23)],data_in[`VWidth*(`APPRam_depth*30+24)-1:`VWidth*(`APPRam_depth*30+23)],data_in[`VWidth*(`APPRam_depth*29+24)-1:`VWidth*(`APPRam_depth*29+23)],data_in[`VWidth*(`APPRam_depth*28+24)-1:`VWidth*(`APPRam_depth*28+23)],data_in[`VWidth*(`APPRam_depth*27+24)-1:`VWidth*(`APPRam_depth*27+23)],data_in[`VWidth*(`APPRam_depth*26+24)-1:`VWidth*(`APPRam_depth*26+23)],data_in[`VWidth*(`APPRam_depth*25+24)-1:`VWidth*(`APPRam_depth*25+23)],data_in[`VWidth*(`APPRam_depth*24+24)-1:`VWidth*(`APPRam_depth*24+23)],data_in[`VWidth*(`APPRam_depth*23+24)-1:`VWidth*(`APPRam_depth*23+23)],data_in[`VWidth*(`APPRam_depth*22+24)-1:`VWidth*(`APPRam_depth*22+23)],data_in[`VWidth*(`APPRam_depth*21+24)-1:`VWidth*(`APPRam_depth*21+23)],data_in[`VWidth*(`APPRam_depth*20+24)-1:`VWidth*(`APPRam_depth*20+23)],data_in[`VWidth*(`APPRam_depth*19+24)-1:`VWidth*(`APPRam_depth*19+23)],data_in[`VWidth*(`APPRam_depth*18+24)-1:`VWidth*(`APPRam_depth*18+23)],data_in[`VWidth*(`APPRam_depth*17+24)-1:`VWidth*(`APPRam_depth*17+23)],data_in[`VWidth*(`APPRam_depth*16+24)-1:`VWidth*(`APPRam_depth*16+23)],data_in[`VWidth*(`APPRam_depth*15+24)-1:`VWidth*(`APPRam_depth*15+23)],data_in[`VWidth*(`APPRam_depth*14+24)-1:`VWidth*(`APPRam_depth*14+23)],data_in[`VWidth*(`APPRam_depth*13+24)-1:`VWidth*(`APPRam_depth*13+23)],data_in[`VWidth*(`APPRam_depth*12+24)-1:`VWidth*(`APPRam_depth*12+23)],data_in[`VWidth*(`APPRam_depth*11+24)-1:`VWidth*(`APPRam_depth*11+23)],data_in[`VWidth*(`APPRam_depth*10+24)-1:`VWidth*(`APPRam_depth*10+23)],data_in[`VWidth*(`APPRam_depth*9+24)-1:`VWidth*(`APPRam_depth*9+23)],data_in[`VWidth*(`APPRam_depth*8+24)-1:`VWidth*(`APPRam_depth*8+23)],data_in[`VWidth*(`APPRam_depth*7+24)-1:`VWidth*(`APPRam_depth*7+23)],data_in[`VWidth*(`APPRam_depth*6+24)-1:`VWidth*(`APPRam_depth*6+23)],data_in[`VWidth*(`APPRam_depth*5+24)-1:`VWidth*(`APPRam_depth*5+23)],data_in[`VWidth*(`APPRam_depth*4+24)-1:`VWidth*(`APPRam_depth*4+23)],data_in[`VWidth*(`APPRam_depth*3+24)-1:`VWidth*(`APPRam_depth*3+23)],data_in[`VWidth*(`APPRam_depth*2+24)-1:`VWidth*(`APPRam_depth*2+23)],data_in[`VWidth*(`APPRam_depth*1+24)-1:`VWidth*(`APPRam_depth*1+23)],data_in[`VWidth*(`APPRam_depth*0+24)-1:`VWidth*(`APPRam_depth*0+23)]};
			end
			24:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+25)-1:`VWidth*(`APPRam_depth*31+24)],data_in[`VWidth*(`APPRam_depth*30+25)-1:`VWidth*(`APPRam_depth*30+24)],data_in[`VWidth*(`APPRam_depth*29+25)-1:`VWidth*(`APPRam_depth*29+24)],data_in[`VWidth*(`APPRam_depth*28+25)-1:`VWidth*(`APPRam_depth*28+24)],data_in[`VWidth*(`APPRam_depth*27+25)-1:`VWidth*(`APPRam_depth*27+24)],data_in[`VWidth*(`APPRam_depth*26+25)-1:`VWidth*(`APPRam_depth*26+24)],data_in[`VWidth*(`APPRam_depth*25+25)-1:`VWidth*(`APPRam_depth*25+24)],data_in[`VWidth*(`APPRam_depth*24+25)-1:`VWidth*(`APPRam_depth*24+24)],data_in[`VWidth*(`APPRam_depth*23+25)-1:`VWidth*(`APPRam_depth*23+24)],data_in[`VWidth*(`APPRam_depth*22+25)-1:`VWidth*(`APPRam_depth*22+24)],data_in[`VWidth*(`APPRam_depth*21+25)-1:`VWidth*(`APPRam_depth*21+24)],data_in[`VWidth*(`APPRam_depth*20+25)-1:`VWidth*(`APPRam_depth*20+24)],data_in[`VWidth*(`APPRam_depth*19+25)-1:`VWidth*(`APPRam_depth*19+24)],data_in[`VWidth*(`APPRam_depth*18+25)-1:`VWidth*(`APPRam_depth*18+24)],data_in[`VWidth*(`APPRam_depth*17+25)-1:`VWidth*(`APPRam_depth*17+24)],data_in[`VWidth*(`APPRam_depth*16+25)-1:`VWidth*(`APPRam_depth*16+24)],data_in[`VWidth*(`APPRam_depth*15+25)-1:`VWidth*(`APPRam_depth*15+24)],data_in[`VWidth*(`APPRam_depth*14+25)-1:`VWidth*(`APPRam_depth*14+24)],data_in[`VWidth*(`APPRam_depth*13+25)-1:`VWidth*(`APPRam_depth*13+24)],data_in[`VWidth*(`APPRam_depth*12+25)-1:`VWidth*(`APPRam_depth*12+24)],data_in[`VWidth*(`APPRam_depth*11+25)-1:`VWidth*(`APPRam_depth*11+24)],data_in[`VWidth*(`APPRam_depth*10+25)-1:`VWidth*(`APPRam_depth*10+24)],data_in[`VWidth*(`APPRam_depth*9+25)-1:`VWidth*(`APPRam_depth*9+24)],data_in[`VWidth*(`APPRam_depth*8+25)-1:`VWidth*(`APPRam_depth*8+24)],data_in[`VWidth*(`APPRam_depth*7+25)-1:`VWidth*(`APPRam_depth*7+24)],data_in[`VWidth*(`APPRam_depth*6+25)-1:`VWidth*(`APPRam_depth*6+24)],data_in[`VWidth*(`APPRam_depth*5+25)-1:`VWidth*(`APPRam_depth*5+24)],data_in[`VWidth*(`APPRam_depth*4+25)-1:`VWidth*(`APPRam_depth*4+24)],data_in[`VWidth*(`APPRam_depth*3+25)-1:`VWidth*(`APPRam_depth*3+24)],data_in[`VWidth*(`APPRam_depth*2+25)-1:`VWidth*(`APPRam_depth*2+24)],data_in[`VWidth*(`APPRam_depth*1+25)-1:`VWidth*(`APPRam_depth*1+24)],data_in[`VWidth*(`APPRam_depth*0+25)-1:`VWidth*(`APPRam_depth*0+24)]};
			end
			25:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+26)-1:`VWidth*(`APPRam_depth*31+25)],data_in[`VWidth*(`APPRam_depth*30+26)-1:`VWidth*(`APPRam_depth*30+25)],data_in[`VWidth*(`APPRam_depth*29+26)-1:`VWidth*(`APPRam_depth*29+25)],data_in[`VWidth*(`APPRam_depth*28+26)-1:`VWidth*(`APPRam_depth*28+25)],data_in[`VWidth*(`APPRam_depth*27+26)-1:`VWidth*(`APPRam_depth*27+25)],data_in[`VWidth*(`APPRam_depth*26+26)-1:`VWidth*(`APPRam_depth*26+25)],data_in[`VWidth*(`APPRam_depth*25+26)-1:`VWidth*(`APPRam_depth*25+25)],data_in[`VWidth*(`APPRam_depth*24+26)-1:`VWidth*(`APPRam_depth*24+25)],data_in[`VWidth*(`APPRam_depth*23+26)-1:`VWidth*(`APPRam_depth*23+25)],data_in[`VWidth*(`APPRam_depth*22+26)-1:`VWidth*(`APPRam_depth*22+25)],data_in[`VWidth*(`APPRam_depth*21+26)-1:`VWidth*(`APPRam_depth*21+25)],data_in[`VWidth*(`APPRam_depth*20+26)-1:`VWidth*(`APPRam_depth*20+25)],data_in[`VWidth*(`APPRam_depth*19+26)-1:`VWidth*(`APPRam_depth*19+25)],data_in[`VWidth*(`APPRam_depth*18+26)-1:`VWidth*(`APPRam_depth*18+25)],data_in[`VWidth*(`APPRam_depth*17+26)-1:`VWidth*(`APPRam_depth*17+25)],data_in[`VWidth*(`APPRam_depth*16+26)-1:`VWidth*(`APPRam_depth*16+25)],data_in[`VWidth*(`APPRam_depth*15+26)-1:`VWidth*(`APPRam_depth*15+25)],data_in[`VWidth*(`APPRam_depth*14+26)-1:`VWidth*(`APPRam_depth*14+25)],data_in[`VWidth*(`APPRam_depth*13+26)-1:`VWidth*(`APPRam_depth*13+25)],data_in[`VWidth*(`APPRam_depth*12+26)-1:`VWidth*(`APPRam_depth*12+25)],data_in[`VWidth*(`APPRam_depth*11+26)-1:`VWidth*(`APPRam_depth*11+25)],data_in[`VWidth*(`APPRam_depth*10+26)-1:`VWidth*(`APPRam_depth*10+25)],data_in[`VWidth*(`APPRam_depth*9+26)-1:`VWidth*(`APPRam_depth*9+25)],data_in[`VWidth*(`APPRam_depth*8+26)-1:`VWidth*(`APPRam_depth*8+25)],data_in[`VWidth*(`APPRam_depth*7+26)-1:`VWidth*(`APPRam_depth*7+25)],data_in[`VWidth*(`APPRam_depth*6+26)-1:`VWidth*(`APPRam_depth*6+25)],data_in[`VWidth*(`APPRam_depth*5+26)-1:`VWidth*(`APPRam_depth*5+25)],data_in[`VWidth*(`APPRam_depth*4+26)-1:`VWidth*(`APPRam_depth*4+25)],data_in[`VWidth*(`APPRam_depth*3+26)-1:`VWidth*(`APPRam_depth*3+25)],data_in[`VWidth*(`APPRam_depth*2+26)-1:`VWidth*(`APPRam_depth*2+25)],data_in[`VWidth*(`APPRam_depth*1+26)-1:`VWidth*(`APPRam_depth*1+25)],data_in[`VWidth*(`APPRam_depth*0+26)-1:`VWidth*(`APPRam_depth*0+25)]};
			end
			26:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+27)-1:`VWidth*(`APPRam_depth*31+26)],data_in[`VWidth*(`APPRam_depth*30+27)-1:`VWidth*(`APPRam_depth*30+26)],data_in[`VWidth*(`APPRam_depth*29+27)-1:`VWidth*(`APPRam_depth*29+26)],data_in[`VWidth*(`APPRam_depth*28+27)-1:`VWidth*(`APPRam_depth*28+26)],data_in[`VWidth*(`APPRam_depth*27+27)-1:`VWidth*(`APPRam_depth*27+26)],data_in[`VWidth*(`APPRam_depth*26+27)-1:`VWidth*(`APPRam_depth*26+26)],data_in[`VWidth*(`APPRam_depth*25+27)-1:`VWidth*(`APPRam_depth*25+26)],data_in[`VWidth*(`APPRam_depth*24+27)-1:`VWidth*(`APPRam_depth*24+26)],data_in[`VWidth*(`APPRam_depth*23+27)-1:`VWidth*(`APPRam_depth*23+26)],data_in[`VWidth*(`APPRam_depth*22+27)-1:`VWidth*(`APPRam_depth*22+26)],data_in[`VWidth*(`APPRam_depth*21+27)-1:`VWidth*(`APPRam_depth*21+26)],data_in[`VWidth*(`APPRam_depth*20+27)-1:`VWidth*(`APPRam_depth*20+26)],data_in[`VWidth*(`APPRam_depth*19+27)-1:`VWidth*(`APPRam_depth*19+26)],data_in[`VWidth*(`APPRam_depth*18+27)-1:`VWidth*(`APPRam_depth*18+26)],data_in[`VWidth*(`APPRam_depth*17+27)-1:`VWidth*(`APPRam_depth*17+26)],data_in[`VWidth*(`APPRam_depth*16+27)-1:`VWidth*(`APPRam_depth*16+26)],data_in[`VWidth*(`APPRam_depth*15+27)-1:`VWidth*(`APPRam_depth*15+26)],data_in[`VWidth*(`APPRam_depth*14+27)-1:`VWidth*(`APPRam_depth*14+26)],data_in[`VWidth*(`APPRam_depth*13+27)-1:`VWidth*(`APPRam_depth*13+26)],data_in[`VWidth*(`APPRam_depth*12+27)-1:`VWidth*(`APPRam_depth*12+26)],data_in[`VWidth*(`APPRam_depth*11+27)-1:`VWidth*(`APPRam_depth*11+26)],data_in[`VWidth*(`APPRam_depth*10+27)-1:`VWidth*(`APPRam_depth*10+26)],data_in[`VWidth*(`APPRam_depth*9+27)-1:`VWidth*(`APPRam_depth*9+26)],data_in[`VWidth*(`APPRam_depth*8+27)-1:`VWidth*(`APPRam_depth*8+26)],data_in[`VWidth*(`APPRam_depth*7+27)-1:`VWidth*(`APPRam_depth*7+26)],data_in[`VWidth*(`APPRam_depth*6+27)-1:`VWidth*(`APPRam_depth*6+26)],data_in[`VWidth*(`APPRam_depth*5+27)-1:`VWidth*(`APPRam_depth*5+26)],data_in[`VWidth*(`APPRam_depth*4+27)-1:`VWidth*(`APPRam_depth*4+26)],data_in[`VWidth*(`APPRam_depth*3+27)-1:`VWidth*(`APPRam_depth*3+26)],data_in[`VWidth*(`APPRam_depth*2+27)-1:`VWidth*(`APPRam_depth*2+26)],data_in[`VWidth*(`APPRam_depth*1+27)-1:`VWidth*(`APPRam_depth*1+26)],data_in[`VWidth*(`APPRam_depth*0+27)-1:`VWidth*(`APPRam_depth*0+26)]};
			end
			27:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+28)-1:`VWidth*(`APPRam_depth*31+27)],data_in[`VWidth*(`APPRam_depth*30+28)-1:`VWidth*(`APPRam_depth*30+27)],data_in[`VWidth*(`APPRam_depth*29+28)-1:`VWidth*(`APPRam_depth*29+27)],data_in[`VWidth*(`APPRam_depth*28+28)-1:`VWidth*(`APPRam_depth*28+27)],data_in[`VWidth*(`APPRam_depth*27+28)-1:`VWidth*(`APPRam_depth*27+27)],data_in[`VWidth*(`APPRam_depth*26+28)-1:`VWidth*(`APPRam_depth*26+27)],data_in[`VWidth*(`APPRam_depth*25+28)-1:`VWidth*(`APPRam_depth*25+27)],data_in[`VWidth*(`APPRam_depth*24+28)-1:`VWidth*(`APPRam_depth*24+27)],data_in[`VWidth*(`APPRam_depth*23+28)-1:`VWidth*(`APPRam_depth*23+27)],data_in[`VWidth*(`APPRam_depth*22+28)-1:`VWidth*(`APPRam_depth*22+27)],data_in[`VWidth*(`APPRam_depth*21+28)-1:`VWidth*(`APPRam_depth*21+27)],data_in[`VWidth*(`APPRam_depth*20+28)-1:`VWidth*(`APPRam_depth*20+27)],data_in[`VWidth*(`APPRam_depth*19+28)-1:`VWidth*(`APPRam_depth*19+27)],data_in[`VWidth*(`APPRam_depth*18+28)-1:`VWidth*(`APPRam_depth*18+27)],data_in[`VWidth*(`APPRam_depth*17+28)-1:`VWidth*(`APPRam_depth*17+27)],data_in[`VWidth*(`APPRam_depth*16+28)-1:`VWidth*(`APPRam_depth*16+27)],data_in[`VWidth*(`APPRam_depth*15+28)-1:`VWidth*(`APPRam_depth*15+27)],data_in[`VWidth*(`APPRam_depth*14+28)-1:`VWidth*(`APPRam_depth*14+27)],data_in[`VWidth*(`APPRam_depth*13+28)-1:`VWidth*(`APPRam_depth*13+27)],data_in[`VWidth*(`APPRam_depth*12+28)-1:`VWidth*(`APPRam_depth*12+27)],data_in[`VWidth*(`APPRam_depth*11+28)-1:`VWidth*(`APPRam_depth*11+27)],data_in[`VWidth*(`APPRam_depth*10+28)-1:`VWidth*(`APPRam_depth*10+27)],data_in[`VWidth*(`APPRam_depth*9+28)-1:`VWidth*(`APPRam_depth*9+27)],data_in[`VWidth*(`APPRam_depth*8+28)-1:`VWidth*(`APPRam_depth*8+27)],data_in[`VWidth*(`APPRam_depth*7+28)-1:`VWidth*(`APPRam_depth*7+27)],data_in[`VWidth*(`APPRam_depth*6+28)-1:`VWidth*(`APPRam_depth*6+27)],data_in[`VWidth*(`APPRam_depth*5+28)-1:`VWidth*(`APPRam_depth*5+27)],data_in[`VWidth*(`APPRam_depth*4+28)-1:`VWidth*(`APPRam_depth*4+27)],data_in[`VWidth*(`APPRam_depth*3+28)-1:`VWidth*(`APPRam_depth*3+27)],data_in[`VWidth*(`APPRam_depth*2+28)-1:`VWidth*(`APPRam_depth*2+27)],data_in[`VWidth*(`APPRam_depth*1+28)-1:`VWidth*(`APPRam_depth*1+27)],data_in[`VWidth*(`APPRam_depth*0+28)-1:`VWidth*(`APPRam_depth*0+27)]};
			end
			28:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+29)-1:`VWidth*(`APPRam_depth*31+28)],data_in[`VWidth*(`APPRam_depth*30+29)-1:`VWidth*(`APPRam_depth*30+28)],data_in[`VWidth*(`APPRam_depth*29+29)-1:`VWidth*(`APPRam_depth*29+28)],data_in[`VWidth*(`APPRam_depth*28+29)-1:`VWidth*(`APPRam_depth*28+28)],data_in[`VWidth*(`APPRam_depth*27+29)-1:`VWidth*(`APPRam_depth*27+28)],data_in[`VWidth*(`APPRam_depth*26+29)-1:`VWidth*(`APPRam_depth*26+28)],data_in[`VWidth*(`APPRam_depth*25+29)-1:`VWidth*(`APPRam_depth*25+28)],data_in[`VWidth*(`APPRam_depth*24+29)-1:`VWidth*(`APPRam_depth*24+28)],data_in[`VWidth*(`APPRam_depth*23+29)-1:`VWidth*(`APPRam_depth*23+28)],data_in[`VWidth*(`APPRam_depth*22+29)-1:`VWidth*(`APPRam_depth*22+28)],data_in[`VWidth*(`APPRam_depth*21+29)-1:`VWidth*(`APPRam_depth*21+28)],data_in[`VWidth*(`APPRam_depth*20+29)-1:`VWidth*(`APPRam_depth*20+28)],data_in[`VWidth*(`APPRam_depth*19+29)-1:`VWidth*(`APPRam_depth*19+28)],data_in[`VWidth*(`APPRam_depth*18+29)-1:`VWidth*(`APPRam_depth*18+28)],data_in[`VWidth*(`APPRam_depth*17+29)-1:`VWidth*(`APPRam_depth*17+28)],data_in[`VWidth*(`APPRam_depth*16+29)-1:`VWidth*(`APPRam_depth*16+28)],data_in[`VWidth*(`APPRam_depth*15+29)-1:`VWidth*(`APPRam_depth*15+28)],data_in[`VWidth*(`APPRam_depth*14+29)-1:`VWidth*(`APPRam_depth*14+28)],data_in[`VWidth*(`APPRam_depth*13+29)-1:`VWidth*(`APPRam_depth*13+28)],data_in[`VWidth*(`APPRam_depth*12+29)-1:`VWidth*(`APPRam_depth*12+28)],data_in[`VWidth*(`APPRam_depth*11+29)-1:`VWidth*(`APPRam_depth*11+28)],data_in[`VWidth*(`APPRam_depth*10+29)-1:`VWidth*(`APPRam_depth*10+28)],data_in[`VWidth*(`APPRam_depth*9+29)-1:`VWidth*(`APPRam_depth*9+28)],data_in[`VWidth*(`APPRam_depth*8+29)-1:`VWidth*(`APPRam_depth*8+28)],data_in[`VWidth*(`APPRam_depth*7+29)-1:`VWidth*(`APPRam_depth*7+28)],data_in[`VWidth*(`APPRam_depth*6+29)-1:`VWidth*(`APPRam_depth*6+28)],data_in[`VWidth*(`APPRam_depth*5+29)-1:`VWidth*(`APPRam_depth*5+28)],data_in[`VWidth*(`APPRam_depth*4+29)-1:`VWidth*(`APPRam_depth*4+28)],data_in[`VWidth*(`APPRam_depth*3+29)-1:`VWidth*(`APPRam_depth*3+28)],data_in[`VWidth*(`APPRam_depth*2+29)-1:`VWidth*(`APPRam_depth*2+28)],data_in[`VWidth*(`APPRam_depth*1+29)-1:`VWidth*(`APPRam_depth*1+28)],data_in[`VWidth*(`APPRam_depth*0+29)-1:`VWidth*(`APPRam_depth*0+28)]};
			end
			29:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+30)-1:`VWidth*(`APPRam_depth*31+29)],data_in[`VWidth*(`APPRam_depth*30+30)-1:`VWidth*(`APPRam_depth*30+29)],data_in[`VWidth*(`APPRam_depth*29+30)-1:`VWidth*(`APPRam_depth*29+29)],data_in[`VWidth*(`APPRam_depth*28+30)-1:`VWidth*(`APPRam_depth*28+29)],data_in[`VWidth*(`APPRam_depth*27+30)-1:`VWidth*(`APPRam_depth*27+29)],data_in[`VWidth*(`APPRam_depth*26+30)-1:`VWidth*(`APPRam_depth*26+29)],data_in[`VWidth*(`APPRam_depth*25+30)-1:`VWidth*(`APPRam_depth*25+29)],data_in[`VWidth*(`APPRam_depth*24+30)-1:`VWidth*(`APPRam_depth*24+29)],data_in[`VWidth*(`APPRam_depth*23+30)-1:`VWidth*(`APPRam_depth*23+29)],data_in[`VWidth*(`APPRam_depth*22+30)-1:`VWidth*(`APPRam_depth*22+29)],data_in[`VWidth*(`APPRam_depth*21+30)-1:`VWidth*(`APPRam_depth*21+29)],data_in[`VWidth*(`APPRam_depth*20+30)-1:`VWidth*(`APPRam_depth*20+29)],data_in[`VWidth*(`APPRam_depth*19+30)-1:`VWidth*(`APPRam_depth*19+29)],data_in[`VWidth*(`APPRam_depth*18+30)-1:`VWidth*(`APPRam_depth*18+29)],data_in[`VWidth*(`APPRam_depth*17+30)-1:`VWidth*(`APPRam_depth*17+29)],data_in[`VWidth*(`APPRam_depth*16+30)-1:`VWidth*(`APPRam_depth*16+29)],data_in[`VWidth*(`APPRam_depth*15+30)-1:`VWidth*(`APPRam_depth*15+29)],data_in[`VWidth*(`APPRam_depth*14+30)-1:`VWidth*(`APPRam_depth*14+29)],data_in[`VWidth*(`APPRam_depth*13+30)-1:`VWidth*(`APPRam_depth*13+29)],data_in[`VWidth*(`APPRam_depth*12+30)-1:`VWidth*(`APPRam_depth*12+29)],data_in[`VWidth*(`APPRam_depth*11+30)-1:`VWidth*(`APPRam_depth*11+29)],data_in[`VWidth*(`APPRam_depth*10+30)-1:`VWidth*(`APPRam_depth*10+29)],data_in[`VWidth*(`APPRam_depth*9+30)-1:`VWidth*(`APPRam_depth*9+29)],data_in[`VWidth*(`APPRam_depth*8+30)-1:`VWidth*(`APPRam_depth*8+29)],data_in[`VWidth*(`APPRam_depth*7+30)-1:`VWidth*(`APPRam_depth*7+29)],data_in[`VWidth*(`APPRam_depth*6+30)-1:`VWidth*(`APPRam_depth*6+29)],data_in[`VWidth*(`APPRam_depth*5+30)-1:`VWidth*(`APPRam_depth*5+29)],data_in[`VWidth*(`APPRam_depth*4+30)-1:`VWidth*(`APPRam_depth*4+29)],data_in[`VWidth*(`APPRam_depth*3+30)-1:`VWidth*(`APPRam_depth*3+29)],data_in[`VWidth*(`APPRam_depth*2+30)-1:`VWidth*(`APPRam_depth*2+29)],data_in[`VWidth*(`APPRam_depth*1+30)-1:`VWidth*(`APPRam_depth*1+29)],data_in[`VWidth*(`APPRam_depth*0+30)-1:`VWidth*(`APPRam_depth*0+29)]};
			end
			30:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+31)-1:`VWidth*(`APPRam_depth*31+30)],data_in[`VWidth*(`APPRam_depth*30+31)-1:`VWidth*(`APPRam_depth*30+30)],data_in[`VWidth*(`APPRam_depth*29+31)-1:`VWidth*(`APPRam_depth*29+30)],data_in[`VWidth*(`APPRam_depth*28+31)-1:`VWidth*(`APPRam_depth*28+30)],data_in[`VWidth*(`APPRam_depth*27+31)-1:`VWidth*(`APPRam_depth*27+30)],data_in[`VWidth*(`APPRam_depth*26+31)-1:`VWidth*(`APPRam_depth*26+30)],data_in[`VWidth*(`APPRam_depth*25+31)-1:`VWidth*(`APPRam_depth*25+30)],data_in[`VWidth*(`APPRam_depth*24+31)-1:`VWidth*(`APPRam_depth*24+30)],data_in[`VWidth*(`APPRam_depth*23+31)-1:`VWidth*(`APPRam_depth*23+30)],data_in[`VWidth*(`APPRam_depth*22+31)-1:`VWidth*(`APPRam_depth*22+30)],data_in[`VWidth*(`APPRam_depth*21+31)-1:`VWidth*(`APPRam_depth*21+30)],data_in[`VWidth*(`APPRam_depth*20+31)-1:`VWidth*(`APPRam_depth*20+30)],data_in[`VWidth*(`APPRam_depth*19+31)-1:`VWidth*(`APPRam_depth*19+30)],data_in[`VWidth*(`APPRam_depth*18+31)-1:`VWidth*(`APPRam_depth*18+30)],data_in[`VWidth*(`APPRam_depth*17+31)-1:`VWidth*(`APPRam_depth*17+30)],data_in[`VWidth*(`APPRam_depth*16+31)-1:`VWidth*(`APPRam_depth*16+30)],data_in[`VWidth*(`APPRam_depth*15+31)-1:`VWidth*(`APPRam_depth*15+30)],data_in[`VWidth*(`APPRam_depth*14+31)-1:`VWidth*(`APPRam_depth*14+30)],data_in[`VWidth*(`APPRam_depth*13+31)-1:`VWidth*(`APPRam_depth*13+30)],data_in[`VWidth*(`APPRam_depth*12+31)-1:`VWidth*(`APPRam_depth*12+30)],data_in[`VWidth*(`APPRam_depth*11+31)-1:`VWidth*(`APPRam_depth*11+30)],data_in[`VWidth*(`APPRam_depth*10+31)-1:`VWidth*(`APPRam_depth*10+30)],data_in[`VWidth*(`APPRam_depth*9+31)-1:`VWidth*(`APPRam_depth*9+30)],data_in[`VWidth*(`APPRam_depth*8+31)-1:`VWidth*(`APPRam_depth*8+30)],data_in[`VWidth*(`APPRam_depth*7+31)-1:`VWidth*(`APPRam_depth*7+30)],data_in[`VWidth*(`APPRam_depth*6+31)-1:`VWidth*(`APPRam_depth*6+30)],data_in[`VWidth*(`APPRam_depth*5+31)-1:`VWidth*(`APPRam_depth*5+30)],data_in[`VWidth*(`APPRam_depth*4+31)-1:`VWidth*(`APPRam_depth*4+30)],data_in[`VWidth*(`APPRam_depth*3+31)-1:`VWidth*(`APPRam_depth*3+30)],data_in[`VWidth*(`APPRam_depth*2+31)-1:`VWidth*(`APPRam_depth*2+30)],data_in[`VWidth*(`APPRam_depth*1+31)-1:`VWidth*(`APPRam_depth*1+30)],data_in[`VWidth*(`APPRam_depth*0+31)-1:`VWidth*(`APPRam_depth*0+30)]};
			end
			31:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+32)-1:`VWidth*(`APPRam_depth*31+31)],data_in[`VWidth*(`APPRam_depth*30+32)-1:`VWidth*(`APPRam_depth*30+31)],data_in[`VWidth*(`APPRam_depth*29+32)-1:`VWidth*(`APPRam_depth*29+31)],data_in[`VWidth*(`APPRam_depth*28+32)-1:`VWidth*(`APPRam_depth*28+31)],data_in[`VWidth*(`APPRam_depth*27+32)-1:`VWidth*(`APPRam_depth*27+31)],data_in[`VWidth*(`APPRam_depth*26+32)-1:`VWidth*(`APPRam_depth*26+31)],data_in[`VWidth*(`APPRam_depth*25+32)-1:`VWidth*(`APPRam_depth*25+31)],data_in[`VWidth*(`APPRam_depth*24+32)-1:`VWidth*(`APPRam_depth*24+31)],data_in[`VWidth*(`APPRam_depth*23+32)-1:`VWidth*(`APPRam_depth*23+31)],data_in[`VWidth*(`APPRam_depth*22+32)-1:`VWidth*(`APPRam_depth*22+31)],data_in[`VWidth*(`APPRam_depth*21+32)-1:`VWidth*(`APPRam_depth*21+31)],data_in[`VWidth*(`APPRam_depth*20+32)-1:`VWidth*(`APPRam_depth*20+31)],data_in[`VWidth*(`APPRam_depth*19+32)-1:`VWidth*(`APPRam_depth*19+31)],data_in[`VWidth*(`APPRam_depth*18+32)-1:`VWidth*(`APPRam_depth*18+31)],data_in[`VWidth*(`APPRam_depth*17+32)-1:`VWidth*(`APPRam_depth*17+31)],data_in[`VWidth*(`APPRam_depth*16+32)-1:`VWidth*(`APPRam_depth*16+31)],data_in[`VWidth*(`APPRam_depth*15+32)-1:`VWidth*(`APPRam_depth*15+31)],data_in[`VWidth*(`APPRam_depth*14+32)-1:`VWidth*(`APPRam_depth*14+31)],data_in[`VWidth*(`APPRam_depth*13+32)-1:`VWidth*(`APPRam_depth*13+31)],data_in[`VWidth*(`APPRam_depth*12+32)-1:`VWidth*(`APPRam_depth*12+31)],data_in[`VWidth*(`APPRam_depth*11+32)-1:`VWidth*(`APPRam_depth*11+31)],data_in[`VWidth*(`APPRam_depth*10+32)-1:`VWidth*(`APPRam_depth*10+31)],data_in[`VWidth*(`APPRam_depth*9+32)-1:`VWidth*(`APPRam_depth*9+31)],data_in[`VWidth*(`APPRam_depth*8+32)-1:`VWidth*(`APPRam_depth*8+31)],data_in[`VWidth*(`APPRam_depth*7+32)-1:`VWidth*(`APPRam_depth*7+31)],data_in[`VWidth*(`APPRam_depth*6+32)-1:`VWidth*(`APPRam_depth*6+31)],data_in[`VWidth*(`APPRam_depth*5+32)-1:`VWidth*(`APPRam_depth*5+31)],data_in[`VWidth*(`APPRam_depth*4+32)-1:`VWidth*(`APPRam_depth*4+31)],data_in[`VWidth*(`APPRam_depth*3+32)-1:`VWidth*(`APPRam_depth*3+31)],data_in[`VWidth*(`APPRam_depth*2+32)-1:`VWidth*(`APPRam_depth*2+31)],data_in[`VWidth*(`APPRam_depth*1+32)-1:`VWidth*(`APPRam_depth*1+31)],data_in[`VWidth*(`APPRam_depth*0+32)-1:`VWidth*(`APPRam_depth*0+31)]};
			end
			32:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+33)-1:`VWidth*(`APPRam_depth*31+32)],data_in[`VWidth*(`APPRam_depth*30+33)-1:`VWidth*(`APPRam_depth*30+32)],data_in[`VWidth*(`APPRam_depth*29+33)-1:`VWidth*(`APPRam_depth*29+32)],data_in[`VWidth*(`APPRam_depth*28+33)-1:`VWidth*(`APPRam_depth*28+32)],data_in[`VWidth*(`APPRam_depth*27+33)-1:`VWidth*(`APPRam_depth*27+32)],data_in[`VWidth*(`APPRam_depth*26+33)-1:`VWidth*(`APPRam_depth*26+32)],data_in[`VWidth*(`APPRam_depth*25+33)-1:`VWidth*(`APPRam_depth*25+32)],data_in[`VWidth*(`APPRam_depth*24+33)-1:`VWidth*(`APPRam_depth*24+32)],data_in[`VWidth*(`APPRam_depth*23+33)-1:`VWidth*(`APPRam_depth*23+32)],data_in[`VWidth*(`APPRam_depth*22+33)-1:`VWidth*(`APPRam_depth*22+32)],data_in[`VWidth*(`APPRam_depth*21+33)-1:`VWidth*(`APPRam_depth*21+32)],data_in[`VWidth*(`APPRam_depth*20+33)-1:`VWidth*(`APPRam_depth*20+32)],data_in[`VWidth*(`APPRam_depth*19+33)-1:`VWidth*(`APPRam_depth*19+32)],data_in[`VWidth*(`APPRam_depth*18+33)-1:`VWidth*(`APPRam_depth*18+32)],data_in[`VWidth*(`APPRam_depth*17+33)-1:`VWidth*(`APPRam_depth*17+32)],data_in[`VWidth*(`APPRam_depth*16+33)-1:`VWidth*(`APPRam_depth*16+32)],data_in[`VWidth*(`APPRam_depth*15+33)-1:`VWidth*(`APPRam_depth*15+32)],data_in[`VWidth*(`APPRam_depth*14+33)-1:`VWidth*(`APPRam_depth*14+32)],data_in[`VWidth*(`APPRam_depth*13+33)-1:`VWidth*(`APPRam_depth*13+32)],data_in[`VWidth*(`APPRam_depth*12+33)-1:`VWidth*(`APPRam_depth*12+32)],data_in[`VWidth*(`APPRam_depth*11+33)-1:`VWidth*(`APPRam_depth*11+32)],data_in[`VWidth*(`APPRam_depth*10+33)-1:`VWidth*(`APPRam_depth*10+32)],data_in[`VWidth*(`APPRam_depth*9+33)-1:`VWidth*(`APPRam_depth*9+32)],data_in[`VWidth*(`APPRam_depth*8+33)-1:`VWidth*(`APPRam_depth*8+32)],data_in[`VWidth*(`APPRam_depth*7+33)-1:`VWidth*(`APPRam_depth*7+32)],data_in[`VWidth*(`APPRam_depth*6+33)-1:`VWidth*(`APPRam_depth*6+32)],data_in[`VWidth*(`APPRam_depth*5+33)-1:`VWidth*(`APPRam_depth*5+32)],data_in[`VWidth*(`APPRam_depth*4+33)-1:`VWidth*(`APPRam_depth*4+32)],data_in[`VWidth*(`APPRam_depth*3+33)-1:`VWidth*(`APPRam_depth*3+32)],data_in[`VWidth*(`APPRam_depth*2+33)-1:`VWidth*(`APPRam_depth*2+32)],data_in[`VWidth*(`APPRam_depth*1+33)-1:`VWidth*(`APPRam_depth*1+32)],data_in[`VWidth*(`APPRam_depth*0+33)-1:`VWidth*(`APPRam_depth*0+32)]};
			end
			33:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+34)-1:`VWidth*(`APPRam_depth*31+33)],data_in[`VWidth*(`APPRam_depth*30+34)-1:`VWidth*(`APPRam_depth*30+33)],data_in[`VWidth*(`APPRam_depth*29+34)-1:`VWidth*(`APPRam_depth*29+33)],data_in[`VWidth*(`APPRam_depth*28+34)-1:`VWidth*(`APPRam_depth*28+33)],data_in[`VWidth*(`APPRam_depth*27+34)-1:`VWidth*(`APPRam_depth*27+33)],data_in[`VWidth*(`APPRam_depth*26+34)-1:`VWidth*(`APPRam_depth*26+33)],data_in[`VWidth*(`APPRam_depth*25+34)-1:`VWidth*(`APPRam_depth*25+33)],data_in[`VWidth*(`APPRam_depth*24+34)-1:`VWidth*(`APPRam_depth*24+33)],data_in[`VWidth*(`APPRam_depth*23+34)-1:`VWidth*(`APPRam_depth*23+33)],data_in[`VWidth*(`APPRam_depth*22+34)-1:`VWidth*(`APPRam_depth*22+33)],data_in[`VWidth*(`APPRam_depth*21+34)-1:`VWidth*(`APPRam_depth*21+33)],data_in[`VWidth*(`APPRam_depth*20+34)-1:`VWidth*(`APPRam_depth*20+33)],data_in[`VWidth*(`APPRam_depth*19+34)-1:`VWidth*(`APPRam_depth*19+33)],data_in[`VWidth*(`APPRam_depth*18+34)-1:`VWidth*(`APPRam_depth*18+33)],data_in[`VWidth*(`APPRam_depth*17+34)-1:`VWidth*(`APPRam_depth*17+33)],data_in[`VWidth*(`APPRam_depth*16+34)-1:`VWidth*(`APPRam_depth*16+33)],data_in[`VWidth*(`APPRam_depth*15+34)-1:`VWidth*(`APPRam_depth*15+33)],data_in[`VWidth*(`APPRam_depth*14+34)-1:`VWidth*(`APPRam_depth*14+33)],data_in[`VWidth*(`APPRam_depth*13+34)-1:`VWidth*(`APPRam_depth*13+33)],data_in[`VWidth*(`APPRam_depth*12+34)-1:`VWidth*(`APPRam_depth*12+33)],data_in[`VWidth*(`APPRam_depth*11+34)-1:`VWidth*(`APPRam_depth*11+33)],data_in[`VWidth*(`APPRam_depth*10+34)-1:`VWidth*(`APPRam_depth*10+33)],data_in[`VWidth*(`APPRam_depth*9+34)-1:`VWidth*(`APPRam_depth*9+33)],data_in[`VWidth*(`APPRam_depth*8+34)-1:`VWidth*(`APPRam_depth*8+33)],data_in[`VWidth*(`APPRam_depth*7+34)-1:`VWidth*(`APPRam_depth*7+33)],data_in[`VWidth*(`APPRam_depth*6+34)-1:`VWidth*(`APPRam_depth*6+33)],data_in[`VWidth*(`APPRam_depth*5+34)-1:`VWidth*(`APPRam_depth*5+33)],data_in[`VWidth*(`APPRam_depth*4+34)-1:`VWidth*(`APPRam_depth*4+33)],data_in[`VWidth*(`APPRam_depth*3+34)-1:`VWidth*(`APPRam_depth*3+33)],data_in[`VWidth*(`APPRam_depth*2+34)-1:`VWidth*(`APPRam_depth*2+33)],data_in[`VWidth*(`APPRam_depth*1+34)-1:`VWidth*(`APPRam_depth*1+33)],data_in[`VWidth*(`APPRam_depth*0+34)-1:`VWidth*(`APPRam_depth*0+33)]};
			end
			34:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+35)-1:`VWidth*(`APPRam_depth*31+34)],data_in[`VWidth*(`APPRam_depth*30+35)-1:`VWidth*(`APPRam_depth*30+34)],data_in[`VWidth*(`APPRam_depth*29+35)-1:`VWidth*(`APPRam_depth*29+34)],data_in[`VWidth*(`APPRam_depth*28+35)-1:`VWidth*(`APPRam_depth*28+34)],data_in[`VWidth*(`APPRam_depth*27+35)-1:`VWidth*(`APPRam_depth*27+34)],data_in[`VWidth*(`APPRam_depth*26+35)-1:`VWidth*(`APPRam_depth*26+34)],data_in[`VWidth*(`APPRam_depth*25+35)-1:`VWidth*(`APPRam_depth*25+34)],data_in[`VWidth*(`APPRam_depth*24+35)-1:`VWidth*(`APPRam_depth*24+34)],data_in[`VWidth*(`APPRam_depth*23+35)-1:`VWidth*(`APPRam_depth*23+34)],data_in[`VWidth*(`APPRam_depth*22+35)-1:`VWidth*(`APPRam_depth*22+34)],data_in[`VWidth*(`APPRam_depth*21+35)-1:`VWidth*(`APPRam_depth*21+34)],data_in[`VWidth*(`APPRam_depth*20+35)-1:`VWidth*(`APPRam_depth*20+34)],data_in[`VWidth*(`APPRam_depth*19+35)-1:`VWidth*(`APPRam_depth*19+34)],data_in[`VWidth*(`APPRam_depth*18+35)-1:`VWidth*(`APPRam_depth*18+34)],data_in[`VWidth*(`APPRam_depth*17+35)-1:`VWidth*(`APPRam_depth*17+34)],data_in[`VWidth*(`APPRam_depth*16+35)-1:`VWidth*(`APPRam_depth*16+34)],data_in[`VWidth*(`APPRam_depth*15+35)-1:`VWidth*(`APPRam_depth*15+34)],data_in[`VWidth*(`APPRam_depth*14+35)-1:`VWidth*(`APPRam_depth*14+34)],data_in[`VWidth*(`APPRam_depth*13+35)-1:`VWidth*(`APPRam_depth*13+34)],data_in[`VWidth*(`APPRam_depth*12+35)-1:`VWidth*(`APPRam_depth*12+34)],data_in[`VWidth*(`APPRam_depth*11+35)-1:`VWidth*(`APPRam_depth*11+34)],data_in[`VWidth*(`APPRam_depth*10+35)-1:`VWidth*(`APPRam_depth*10+34)],data_in[`VWidth*(`APPRam_depth*9+35)-1:`VWidth*(`APPRam_depth*9+34)],data_in[`VWidth*(`APPRam_depth*8+35)-1:`VWidth*(`APPRam_depth*8+34)],data_in[`VWidth*(`APPRam_depth*7+35)-1:`VWidth*(`APPRam_depth*7+34)],data_in[`VWidth*(`APPRam_depth*6+35)-1:`VWidth*(`APPRam_depth*6+34)],data_in[`VWidth*(`APPRam_depth*5+35)-1:`VWidth*(`APPRam_depth*5+34)],data_in[`VWidth*(`APPRam_depth*4+35)-1:`VWidth*(`APPRam_depth*4+34)],data_in[`VWidth*(`APPRam_depth*3+35)-1:`VWidth*(`APPRam_depth*3+34)],data_in[`VWidth*(`APPRam_depth*2+35)-1:`VWidth*(`APPRam_depth*2+34)],data_in[`VWidth*(`APPRam_depth*1+35)-1:`VWidth*(`APPRam_depth*1+34)],data_in[`VWidth*(`APPRam_depth*0+35)-1:`VWidth*(`APPRam_depth*0+34)]};
			end
			35:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+36)-1:`VWidth*(`APPRam_depth*31+35)],data_in[`VWidth*(`APPRam_depth*30+36)-1:`VWidth*(`APPRam_depth*30+35)],data_in[`VWidth*(`APPRam_depth*29+36)-1:`VWidth*(`APPRam_depth*29+35)],data_in[`VWidth*(`APPRam_depth*28+36)-1:`VWidth*(`APPRam_depth*28+35)],data_in[`VWidth*(`APPRam_depth*27+36)-1:`VWidth*(`APPRam_depth*27+35)],data_in[`VWidth*(`APPRam_depth*26+36)-1:`VWidth*(`APPRam_depth*26+35)],data_in[`VWidth*(`APPRam_depth*25+36)-1:`VWidth*(`APPRam_depth*25+35)],data_in[`VWidth*(`APPRam_depth*24+36)-1:`VWidth*(`APPRam_depth*24+35)],data_in[`VWidth*(`APPRam_depth*23+36)-1:`VWidth*(`APPRam_depth*23+35)],data_in[`VWidth*(`APPRam_depth*22+36)-1:`VWidth*(`APPRam_depth*22+35)],data_in[`VWidth*(`APPRam_depth*21+36)-1:`VWidth*(`APPRam_depth*21+35)],data_in[`VWidth*(`APPRam_depth*20+36)-1:`VWidth*(`APPRam_depth*20+35)],data_in[`VWidth*(`APPRam_depth*19+36)-1:`VWidth*(`APPRam_depth*19+35)],data_in[`VWidth*(`APPRam_depth*18+36)-1:`VWidth*(`APPRam_depth*18+35)],data_in[`VWidth*(`APPRam_depth*17+36)-1:`VWidth*(`APPRam_depth*17+35)],data_in[`VWidth*(`APPRam_depth*16+36)-1:`VWidth*(`APPRam_depth*16+35)],data_in[`VWidth*(`APPRam_depth*15+36)-1:`VWidth*(`APPRam_depth*15+35)],data_in[`VWidth*(`APPRam_depth*14+36)-1:`VWidth*(`APPRam_depth*14+35)],data_in[`VWidth*(`APPRam_depth*13+36)-1:`VWidth*(`APPRam_depth*13+35)],data_in[`VWidth*(`APPRam_depth*12+36)-1:`VWidth*(`APPRam_depth*12+35)],data_in[`VWidth*(`APPRam_depth*11+36)-1:`VWidth*(`APPRam_depth*11+35)],data_in[`VWidth*(`APPRam_depth*10+36)-1:`VWidth*(`APPRam_depth*10+35)],data_in[`VWidth*(`APPRam_depth*9+36)-1:`VWidth*(`APPRam_depth*9+35)],data_in[`VWidth*(`APPRam_depth*8+36)-1:`VWidth*(`APPRam_depth*8+35)],data_in[`VWidth*(`APPRam_depth*7+36)-1:`VWidth*(`APPRam_depth*7+35)],data_in[`VWidth*(`APPRam_depth*6+36)-1:`VWidth*(`APPRam_depth*6+35)],data_in[`VWidth*(`APPRam_depth*5+36)-1:`VWidth*(`APPRam_depth*5+35)],data_in[`VWidth*(`APPRam_depth*4+36)-1:`VWidth*(`APPRam_depth*4+35)],data_in[`VWidth*(`APPRam_depth*3+36)-1:`VWidth*(`APPRam_depth*3+35)],data_in[`VWidth*(`APPRam_depth*2+36)-1:`VWidth*(`APPRam_depth*2+35)],data_in[`VWidth*(`APPRam_depth*1+36)-1:`VWidth*(`APPRam_depth*1+35)],data_in[`VWidth*(`APPRam_depth*0+36)-1:`VWidth*(`APPRam_depth*0+35)]};
			end
			36:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+37)-1:`VWidth*(`APPRam_depth*31+36)],data_in[`VWidth*(`APPRam_depth*30+37)-1:`VWidth*(`APPRam_depth*30+36)],data_in[`VWidth*(`APPRam_depth*29+37)-1:`VWidth*(`APPRam_depth*29+36)],data_in[`VWidth*(`APPRam_depth*28+37)-1:`VWidth*(`APPRam_depth*28+36)],data_in[`VWidth*(`APPRam_depth*27+37)-1:`VWidth*(`APPRam_depth*27+36)],data_in[`VWidth*(`APPRam_depth*26+37)-1:`VWidth*(`APPRam_depth*26+36)],data_in[`VWidth*(`APPRam_depth*25+37)-1:`VWidth*(`APPRam_depth*25+36)],data_in[`VWidth*(`APPRam_depth*24+37)-1:`VWidth*(`APPRam_depth*24+36)],data_in[`VWidth*(`APPRam_depth*23+37)-1:`VWidth*(`APPRam_depth*23+36)],data_in[`VWidth*(`APPRam_depth*22+37)-1:`VWidth*(`APPRam_depth*22+36)],data_in[`VWidth*(`APPRam_depth*21+37)-1:`VWidth*(`APPRam_depth*21+36)],data_in[`VWidth*(`APPRam_depth*20+37)-1:`VWidth*(`APPRam_depth*20+36)],data_in[`VWidth*(`APPRam_depth*19+37)-1:`VWidth*(`APPRam_depth*19+36)],data_in[`VWidth*(`APPRam_depth*18+37)-1:`VWidth*(`APPRam_depth*18+36)],data_in[`VWidth*(`APPRam_depth*17+37)-1:`VWidth*(`APPRam_depth*17+36)],data_in[`VWidth*(`APPRam_depth*16+37)-1:`VWidth*(`APPRam_depth*16+36)],data_in[`VWidth*(`APPRam_depth*15+37)-1:`VWidth*(`APPRam_depth*15+36)],data_in[`VWidth*(`APPRam_depth*14+37)-1:`VWidth*(`APPRam_depth*14+36)],data_in[`VWidth*(`APPRam_depth*13+37)-1:`VWidth*(`APPRam_depth*13+36)],data_in[`VWidth*(`APPRam_depth*12+37)-1:`VWidth*(`APPRam_depth*12+36)],data_in[`VWidth*(`APPRam_depth*11+37)-1:`VWidth*(`APPRam_depth*11+36)],data_in[`VWidth*(`APPRam_depth*10+37)-1:`VWidth*(`APPRam_depth*10+36)],data_in[`VWidth*(`APPRam_depth*9+37)-1:`VWidth*(`APPRam_depth*9+36)],data_in[`VWidth*(`APPRam_depth*8+37)-1:`VWidth*(`APPRam_depth*8+36)],data_in[`VWidth*(`APPRam_depth*7+37)-1:`VWidth*(`APPRam_depth*7+36)],data_in[`VWidth*(`APPRam_depth*6+37)-1:`VWidth*(`APPRam_depth*6+36)],data_in[`VWidth*(`APPRam_depth*5+37)-1:`VWidth*(`APPRam_depth*5+36)],data_in[`VWidth*(`APPRam_depth*4+37)-1:`VWidth*(`APPRam_depth*4+36)],data_in[`VWidth*(`APPRam_depth*3+37)-1:`VWidth*(`APPRam_depth*3+36)],data_in[`VWidth*(`APPRam_depth*2+37)-1:`VWidth*(`APPRam_depth*2+36)],data_in[`VWidth*(`APPRam_depth*1+37)-1:`VWidth*(`APPRam_depth*1+36)],data_in[`VWidth*(`APPRam_depth*0+37)-1:`VWidth*(`APPRam_depth*0+36)]};
			end
			37:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+38)-1:`VWidth*(`APPRam_depth*31+37)],data_in[`VWidth*(`APPRam_depth*30+38)-1:`VWidth*(`APPRam_depth*30+37)],data_in[`VWidth*(`APPRam_depth*29+38)-1:`VWidth*(`APPRam_depth*29+37)],data_in[`VWidth*(`APPRam_depth*28+38)-1:`VWidth*(`APPRam_depth*28+37)],data_in[`VWidth*(`APPRam_depth*27+38)-1:`VWidth*(`APPRam_depth*27+37)],data_in[`VWidth*(`APPRam_depth*26+38)-1:`VWidth*(`APPRam_depth*26+37)],data_in[`VWidth*(`APPRam_depth*25+38)-1:`VWidth*(`APPRam_depth*25+37)],data_in[`VWidth*(`APPRam_depth*24+38)-1:`VWidth*(`APPRam_depth*24+37)],data_in[`VWidth*(`APPRam_depth*23+38)-1:`VWidth*(`APPRam_depth*23+37)],data_in[`VWidth*(`APPRam_depth*22+38)-1:`VWidth*(`APPRam_depth*22+37)],data_in[`VWidth*(`APPRam_depth*21+38)-1:`VWidth*(`APPRam_depth*21+37)],data_in[`VWidth*(`APPRam_depth*20+38)-1:`VWidth*(`APPRam_depth*20+37)],data_in[`VWidth*(`APPRam_depth*19+38)-1:`VWidth*(`APPRam_depth*19+37)],data_in[`VWidth*(`APPRam_depth*18+38)-1:`VWidth*(`APPRam_depth*18+37)],data_in[`VWidth*(`APPRam_depth*17+38)-1:`VWidth*(`APPRam_depth*17+37)],data_in[`VWidth*(`APPRam_depth*16+38)-1:`VWidth*(`APPRam_depth*16+37)],data_in[`VWidth*(`APPRam_depth*15+38)-1:`VWidth*(`APPRam_depth*15+37)],data_in[`VWidth*(`APPRam_depth*14+38)-1:`VWidth*(`APPRam_depth*14+37)],data_in[`VWidth*(`APPRam_depth*13+38)-1:`VWidth*(`APPRam_depth*13+37)],data_in[`VWidth*(`APPRam_depth*12+38)-1:`VWidth*(`APPRam_depth*12+37)],data_in[`VWidth*(`APPRam_depth*11+38)-1:`VWidth*(`APPRam_depth*11+37)],data_in[`VWidth*(`APPRam_depth*10+38)-1:`VWidth*(`APPRam_depth*10+37)],data_in[`VWidth*(`APPRam_depth*9+38)-1:`VWidth*(`APPRam_depth*9+37)],data_in[`VWidth*(`APPRam_depth*8+38)-1:`VWidth*(`APPRam_depth*8+37)],data_in[`VWidth*(`APPRam_depth*7+38)-1:`VWidth*(`APPRam_depth*7+37)],data_in[`VWidth*(`APPRam_depth*6+38)-1:`VWidth*(`APPRam_depth*6+37)],data_in[`VWidth*(`APPRam_depth*5+38)-1:`VWidth*(`APPRam_depth*5+37)],data_in[`VWidth*(`APPRam_depth*4+38)-1:`VWidth*(`APPRam_depth*4+37)],data_in[`VWidth*(`APPRam_depth*3+38)-1:`VWidth*(`APPRam_depth*3+37)],data_in[`VWidth*(`APPRam_depth*2+38)-1:`VWidth*(`APPRam_depth*2+37)],data_in[`VWidth*(`APPRam_depth*1+38)-1:`VWidth*(`APPRam_depth*1+37)],data_in[`VWidth*(`APPRam_depth*0+38)-1:`VWidth*(`APPRam_depth*0+37)]};
			end
			38:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+39)-1:`VWidth*(`APPRam_depth*31+38)],data_in[`VWidth*(`APPRam_depth*30+39)-1:`VWidth*(`APPRam_depth*30+38)],data_in[`VWidth*(`APPRam_depth*29+39)-1:`VWidth*(`APPRam_depth*29+38)],data_in[`VWidth*(`APPRam_depth*28+39)-1:`VWidth*(`APPRam_depth*28+38)],data_in[`VWidth*(`APPRam_depth*27+39)-1:`VWidth*(`APPRam_depth*27+38)],data_in[`VWidth*(`APPRam_depth*26+39)-1:`VWidth*(`APPRam_depth*26+38)],data_in[`VWidth*(`APPRam_depth*25+39)-1:`VWidth*(`APPRam_depth*25+38)],data_in[`VWidth*(`APPRam_depth*24+39)-1:`VWidth*(`APPRam_depth*24+38)],data_in[`VWidth*(`APPRam_depth*23+39)-1:`VWidth*(`APPRam_depth*23+38)],data_in[`VWidth*(`APPRam_depth*22+39)-1:`VWidth*(`APPRam_depth*22+38)],data_in[`VWidth*(`APPRam_depth*21+39)-1:`VWidth*(`APPRam_depth*21+38)],data_in[`VWidth*(`APPRam_depth*20+39)-1:`VWidth*(`APPRam_depth*20+38)],data_in[`VWidth*(`APPRam_depth*19+39)-1:`VWidth*(`APPRam_depth*19+38)],data_in[`VWidth*(`APPRam_depth*18+39)-1:`VWidth*(`APPRam_depth*18+38)],data_in[`VWidth*(`APPRam_depth*17+39)-1:`VWidth*(`APPRam_depth*17+38)],data_in[`VWidth*(`APPRam_depth*16+39)-1:`VWidth*(`APPRam_depth*16+38)],data_in[`VWidth*(`APPRam_depth*15+39)-1:`VWidth*(`APPRam_depth*15+38)],data_in[`VWidth*(`APPRam_depth*14+39)-1:`VWidth*(`APPRam_depth*14+38)],data_in[`VWidth*(`APPRam_depth*13+39)-1:`VWidth*(`APPRam_depth*13+38)],data_in[`VWidth*(`APPRam_depth*12+39)-1:`VWidth*(`APPRam_depth*12+38)],data_in[`VWidth*(`APPRam_depth*11+39)-1:`VWidth*(`APPRam_depth*11+38)],data_in[`VWidth*(`APPRam_depth*10+39)-1:`VWidth*(`APPRam_depth*10+38)],data_in[`VWidth*(`APPRam_depth*9+39)-1:`VWidth*(`APPRam_depth*9+38)],data_in[`VWidth*(`APPRam_depth*8+39)-1:`VWidth*(`APPRam_depth*8+38)],data_in[`VWidth*(`APPRam_depth*7+39)-1:`VWidth*(`APPRam_depth*7+38)],data_in[`VWidth*(`APPRam_depth*6+39)-1:`VWidth*(`APPRam_depth*6+38)],data_in[`VWidth*(`APPRam_depth*5+39)-1:`VWidth*(`APPRam_depth*5+38)],data_in[`VWidth*(`APPRam_depth*4+39)-1:`VWidth*(`APPRam_depth*4+38)],data_in[`VWidth*(`APPRam_depth*3+39)-1:`VWidth*(`APPRam_depth*3+38)],data_in[`VWidth*(`APPRam_depth*2+39)-1:`VWidth*(`APPRam_depth*2+38)],data_in[`VWidth*(`APPRam_depth*1+39)-1:`VWidth*(`APPRam_depth*1+38)],data_in[`VWidth*(`APPRam_depth*0+39)-1:`VWidth*(`APPRam_depth*0+38)]};
			end
			39:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+40)-1:`VWidth*(`APPRam_depth*31+39)],data_in[`VWidth*(`APPRam_depth*30+40)-1:`VWidth*(`APPRam_depth*30+39)],data_in[`VWidth*(`APPRam_depth*29+40)-1:`VWidth*(`APPRam_depth*29+39)],data_in[`VWidth*(`APPRam_depth*28+40)-1:`VWidth*(`APPRam_depth*28+39)],data_in[`VWidth*(`APPRam_depth*27+40)-1:`VWidth*(`APPRam_depth*27+39)],data_in[`VWidth*(`APPRam_depth*26+40)-1:`VWidth*(`APPRam_depth*26+39)],data_in[`VWidth*(`APPRam_depth*25+40)-1:`VWidth*(`APPRam_depth*25+39)],data_in[`VWidth*(`APPRam_depth*24+40)-1:`VWidth*(`APPRam_depth*24+39)],data_in[`VWidth*(`APPRam_depth*23+40)-1:`VWidth*(`APPRam_depth*23+39)],data_in[`VWidth*(`APPRam_depth*22+40)-1:`VWidth*(`APPRam_depth*22+39)],data_in[`VWidth*(`APPRam_depth*21+40)-1:`VWidth*(`APPRam_depth*21+39)],data_in[`VWidth*(`APPRam_depth*20+40)-1:`VWidth*(`APPRam_depth*20+39)],data_in[`VWidth*(`APPRam_depth*19+40)-1:`VWidth*(`APPRam_depth*19+39)],data_in[`VWidth*(`APPRam_depth*18+40)-1:`VWidth*(`APPRam_depth*18+39)],data_in[`VWidth*(`APPRam_depth*17+40)-1:`VWidth*(`APPRam_depth*17+39)],data_in[`VWidth*(`APPRam_depth*16+40)-1:`VWidth*(`APPRam_depth*16+39)],data_in[`VWidth*(`APPRam_depth*15+40)-1:`VWidth*(`APPRam_depth*15+39)],data_in[`VWidth*(`APPRam_depth*14+40)-1:`VWidth*(`APPRam_depth*14+39)],data_in[`VWidth*(`APPRam_depth*13+40)-1:`VWidth*(`APPRam_depth*13+39)],data_in[`VWidth*(`APPRam_depth*12+40)-1:`VWidth*(`APPRam_depth*12+39)],data_in[`VWidth*(`APPRam_depth*11+40)-1:`VWidth*(`APPRam_depth*11+39)],data_in[`VWidth*(`APPRam_depth*10+40)-1:`VWidth*(`APPRam_depth*10+39)],data_in[`VWidth*(`APPRam_depth*9+40)-1:`VWidth*(`APPRam_depth*9+39)],data_in[`VWidth*(`APPRam_depth*8+40)-1:`VWidth*(`APPRam_depth*8+39)],data_in[`VWidth*(`APPRam_depth*7+40)-1:`VWidth*(`APPRam_depth*7+39)],data_in[`VWidth*(`APPRam_depth*6+40)-1:`VWidth*(`APPRam_depth*6+39)],data_in[`VWidth*(`APPRam_depth*5+40)-1:`VWidth*(`APPRam_depth*5+39)],data_in[`VWidth*(`APPRam_depth*4+40)-1:`VWidth*(`APPRam_depth*4+39)],data_in[`VWidth*(`APPRam_depth*3+40)-1:`VWidth*(`APPRam_depth*3+39)],data_in[`VWidth*(`APPRam_depth*2+40)-1:`VWidth*(`APPRam_depth*2+39)],data_in[`VWidth*(`APPRam_depth*1+40)-1:`VWidth*(`APPRam_depth*1+39)],data_in[`VWidth*(`APPRam_depth*0+40)-1:`VWidth*(`APPRam_depth*0+39)]};
			end
			40:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+41)-1:`VWidth*(`APPRam_depth*31+40)],data_in[`VWidth*(`APPRam_depth*30+41)-1:`VWidth*(`APPRam_depth*30+40)],data_in[`VWidth*(`APPRam_depth*29+41)-1:`VWidth*(`APPRam_depth*29+40)],data_in[`VWidth*(`APPRam_depth*28+41)-1:`VWidth*(`APPRam_depth*28+40)],data_in[`VWidth*(`APPRam_depth*27+41)-1:`VWidth*(`APPRam_depth*27+40)],data_in[`VWidth*(`APPRam_depth*26+41)-1:`VWidth*(`APPRam_depth*26+40)],data_in[`VWidth*(`APPRam_depth*25+41)-1:`VWidth*(`APPRam_depth*25+40)],data_in[`VWidth*(`APPRam_depth*24+41)-1:`VWidth*(`APPRam_depth*24+40)],data_in[`VWidth*(`APPRam_depth*23+41)-1:`VWidth*(`APPRam_depth*23+40)],data_in[`VWidth*(`APPRam_depth*22+41)-1:`VWidth*(`APPRam_depth*22+40)],data_in[`VWidth*(`APPRam_depth*21+41)-1:`VWidth*(`APPRam_depth*21+40)],data_in[`VWidth*(`APPRam_depth*20+41)-1:`VWidth*(`APPRam_depth*20+40)],data_in[`VWidth*(`APPRam_depth*19+41)-1:`VWidth*(`APPRam_depth*19+40)],data_in[`VWidth*(`APPRam_depth*18+41)-1:`VWidth*(`APPRam_depth*18+40)],data_in[`VWidth*(`APPRam_depth*17+41)-1:`VWidth*(`APPRam_depth*17+40)],data_in[`VWidth*(`APPRam_depth*16+41)-1:`VWidth*(`APPRam_depth*16+40)],data_in[`VWidth*(`APPRam_depth*15+41)-1:`VWidth*(`APPRam_depth*15+40)],data_in[`VWidth*(`APPRam_depth*14+41)-1:`VWidth*(`APPRam_depth*14+40)],data_in[`VWidth*(`APPRam_depth*13+41)-1:`VWidth*(`APPRam_depth*13+40)],data_in[`VWidth*(`APPRam_depth*12+41)-1:`VWidth*(`APPRam_depth*12+40)],data_in[`VWidth*(`APPRam_depth*11+41)-1:`VWidth*(`APPRam_depth*11+40)],data_in[`VWidth*(`APPRam_depth*10+41)-1:`VWidth*(`APPRam_depth*10+40)],data_in[`VWidth*(`APPRam_depth*9+41)-1:`VWidth*(`APPRam_depth*9+40)],data_in[`VWidth*(`APPRam_depth*8+41)-1:`VWidth*(`APPRam_depth*8+40)],data_in[`VWidth*(`APPRam_depth*7+41)-1:`VWidth*(`APPRam_depth*7+40)],data_in[`VWidth*(`APPRam_depth*6+41)-1:`VWidth*(`APPRam_depth*6+40)],data_in[`VWidth*(`APPRam_depth*5+41)-1:`VWidth*(`APPRam_depth*5+40)],data_in[`VWidth*(`APPRam_depth*4+41)-1:`VWidth*(`APPRam_depth*4+40)],data_in[`VWidth*(`APPRam_depth*3+41)-1:`VWidth*(`APPRam_depth*3+40)],data_in[`VWidth*(`APPRam_depth*2+41)-1:`VWidth*(`APPRam_depth*2+40)],data_in[`VWidth*(`APPRam_depth*1+41)-1:`VWidth*(`APPRam_depth*1+40)],data_in[`VWidth*(`APPRam_depth*0+41)-1:`VWidth*(`APPRam_depth*0+40)]};
			end
			41:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+42)-1:`VWidth*(`APPRam_depth*31+41)],data_in[`VWidth*(`APPRam_depth*30+42)-1:`VWidth*(`APPRam_depth*30+41)],data_in[`VWidth*(`APPRam_depth*29+42)-1:`VWidth*(`APPRam_depth*29+41)],data_in[`VWidth*(`APPRam_depth*28+42)-1:`VWidth*(`APPRam_depth*28+41)],data_in[`VWidth*(`APPRam_depth*27+42)-1:`VWidth*(`APPRam_depth*27+41)],data_in[`VWidth*(`APPRam_depth*26+42)-1:`VWidth*(`APPRam_depth*26+41)],data_in[`VWidth*(`APPRam_depth*25+42)-1:`VWidth*(`APPRam_depth*25+41)],data_in[`VWidth*(`APPRam_depth*24+42)-1:`VWidth*(`APPRam_depth*24+41)],data_in[`VWidth*(`APPRam_depth*23+42)-1:`VWidth*(`APPRam_depth*23+41)],data_in[`VWidth*(`APPRam_depth*22+42)-1:`VWidth*(`APPRam_depth*22+41)],data_in[`VWidth*(`APPRam_depth*21+42)-1:`VWidth*(`APPRam_depth*21+41)],data_in[`VWidth*(`APPRam_depth*20+42)-1:`VWidth*(`APPRam_depth*20+41)],data_in[`VWidth*(`APPRam_depth*19+42)-1:`VWidth*(`APPRam_depth*19+41)],data_in[`VWidth*(`APPRam_depth*18+42)-1:`VWidth*(`APPRam_depth*18+41)],data_in[`VWidth*(`APPRam_depth*17+42)-1:`VWidth*(`APPRam_depth*17+41)],data_in[`VWidth*(`APPRam_depth*16+42)-1:`VWidth*(`APPRam_depth*16+41)],data_in[`VWidth*(`APPRam_depth*15+42)-1:`VWidth*(`APPRam_depth*15+41)],data_in[`VWidth*(`APPRam_depth*14+42)-1:`VWidth*(`APPRam_depth*14+41)],data_in[`VWidth*(`APPRam_depth*13+42)-1:`VWidth*(`APPRam_depth*13+41)],data_in[`VWidth*(`APPRam_depth*12+42)-1:`VWidth*(`APPRam_depth*12+41)],data_in[`VWidth*(`APPRam_depth*11+42)-1:`VWidth*(`APPRam_depth*11+41)],data_in[`VWidth*(`APPRam_depth*10+42)-1:`VWidth*(`APPRam_depth*10+41)],data_in[`VWidth*(`APPRam_depth*9+42)-1:`VWidth*(`APPRam_depth*9+41)],data_in[`VWidth*(`APPRam_depth*8+42)-1:`VWidth*(`APPRam_depth*8+41)],data_in[`VWidth*(`APPRam_depth*7+42)-1:`VWidth*(`APPRam_depth*7+41)],data_in[`VWidth*(`APPRam_depth*6+42)-1:`VWidth*(`APPRam_depth*6+41)],data_in[`VWidth*(`APPRam_depth*5+42)-1:`VWidth*(`APPRam_depth*5+41)],data_in[`VWidth*(`APPRam_depth*4+42)-1:`VWidth*(`APPRam_depth*4+41)],data_in[`VWidth*(`APPRam_depth*3+42)-1:`VWidth*(`APPRam_depth*3+41)],data_in[`VWidth*(`APPRam_depth*2+42)-1:`VWidth*(`APPRam_depth*2+41)],data_in[`VWidth*(`APPRam_depth*1+42)-1:`VWidth*(`APPRam_depth*1+41)],data_in[`VWidth*(`APPRam_depth*0+42)-1:`VWidth*(`APPRam_depth*0+41)]};
			end
			42:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+43)-1:`VWidth*(`APPRam_depth*31+42)],data_in[`VWidth*(`APPRam_depth*30+43)-1:`VWidth*(`APPRam_depth*30+42)],data_in[`VWidth*(`APPRam_depth*29+43)-1:`VWidth*(`APPRam_depth*29+42)],data_in[`VWidth*(`APPRam_depth*28+43)-1:`VWidth*(`APPRam_depth*28+42)],data_in[`VWidth*(`APPRam_depth*27+43)-1:`VWidth*(`APPRam_depth*27+42)],data_in[`VWidth*(`APPRam_depth*26+43)-1:`VWidth*(`APPRam_depth*26+42)],data_in[`VWidth*(`APPRam_depth*25+43)-1:`VWidth*(`APPRam_depth*25+42)],data_in[`VWidth*(`APPRam_depth*24+43)-1:`VWidth*(`APPRam_depth*24+42)],data_in[`VWidth*(`APPRam_depth*23+43)-1:`VWidth*(`APPRam_depth*23+42)],data_in[`VWidth*(`APPRam_depth*22+43)-1:`VWidth*(`APPRam_depth*22+42)],data_in[`VWidth*(`APPRam_depth*21+43)-1:`VWidth*(`APPRam_depth*21+42)],data_in[`VWidth*(`APPRam_depth*20+43)-1:`VWidth*(`APPRam_depth*20+42)],data_in[`VWidth*(`APPRam_depth*19+43)-1:`VWidth*(`APPRam_depth*19+42)],data_in[`VWidth*(`APPRam_depth*18+43)-1:`VWidth*(`APPRam_depth*18+42)],data_in[`VWidth*(`APPRam_depth*17+43)-1:`VWidth*(`APPRam_depth*17+42)],data_in[`VWidth*(`APPRam_depth*16+43)-1:`VWidth*(`APPRam_depth*16+42)],data_in[`VWidth*(`APPRam_depth*15+43)-1:`VWidth*(`APPRam_depth*15+42)],data_in[`VWidth*(`APPRam_depth*14+43)-1:`VWidth*(`APPRam_depth*14+42)],data_in[`VWidth*(`APPRam_depth*13+43)-1:`VWidth*(`APPRam_depth*13+42)],data_in[`VWidth*(`APPRam_depth*12+43)-1:`VWidth*(`APPRam_depth*12+42)],data_in[`VWidth*(`APPRam_depth*11+43)-1:`VWidth*(`APPRam_depth*11+42)],data_in[`VWidth*(`APPRam_depth*10+43)-1:`VWidth*(`APPRam_depth*10+42)],data_in[`VWidth*(`APPRam_depth*9+43)-1:`VWidth*(`APPRam_depth*9+42)],data_in[`VWidth*(`APPRam_depth*8+43)-1:`VWidth*(`APPRam_depth*8+42)],data_in[`VWidth*(`APPRam_depth*7+43)-1:`VWidth*(`APPRam_depth*7+42)],data_in[`VWidth*(`APPRam_depth*6+43)-1:`VWidth*(`APPRam_depth*6+42)],data_in[`VWidth*(`APPRam_depth*5+43)-1:`VWidth*(`APPRam_depth*5+42)],data_in[`VWidth*(`APPRam_depth*4+43)-1:`VWidth*(`APPRam_depth*4+42)],data_in[`VWidth*(`APPRam_depth*3+43)-1:`VWidth*(`APPRam_depth*3+42)],data_in[`VWidth*(`APPRam_depth*2+43)-1:`VWidth*(`APPRam_depth*2+42)],data_in[`VWidth*(`APPRam_depth*1+43)-1:`VWidth*(`APPRam_depth*1+42)],data_in[`VWidth*(`APPRam_depth*0+43)-1:`VWidth*(`APPRam_depth*0+42)]};
			end
			43:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+44)-1:`VWidth*(`APPRam_depth*31+43)],data_in[`VWidth*(`APPRam_depth*30+44)-1:`VWidth*(`APPRam_depth*30+43)],data_in[`VWidth*(`APPRam_depth*29+44)-1:`VWidth*(`APPRam_depth*29+43)],data_in[`VWidth*(`APPRam_depth*28+44)-1:`VWidth*(`APPRam_depth*28+43)],data_in[`VWidth*(`APPRam_depth*27+44)-1:`VWidth*(`APPRam_depth*27+43)],data_in[`VWidth*(`APPRam_depth*26+44)-1:`VWidth*(`APPRam_depth*26+43)],data_in[`VWidth*(`APPRam_depth*25+44)-1:`VWidth*(`APPRam_depth*25+43)],data_in[`VWidth*(`APPRam_depth*24+44)-1:`VWidth*(`APPRam_depth*24+43)],data_in[`VWidth*(`APPRam_depth*23+44)-1:`VWidth*(`APPRam_depth*23+43)],data_in[`VWidth*(`APPRam_depth*22+44)-1:`VWidth*(`APPRam_depth*22+43)],data_in[`VWidth*(`APPRam_depth*21+44)-1:`VWidth*(`APPRam_depth*21+43)],data_in[`VWidth*(`APPRam_depth*20+44)-1:`VWidth*(`APPRam_depth*20+43)],data_in[`VWidth*(`APPRam_depth*19+44)-1:`VWidth*(`APPRam_depth*19+43)],data_in[`VWidth*(`APPRam_depth*18+44)-1:`VWidth*(`APPRam_depth*18+43)],data_in[`VWidth*(`APPRam_depth*17+44)-1:`VWidth*(`APPRam_depth*17+43)],data_in[`VWidth*(`APPRam_depth*16+44)-1:`VWidth*(`APPRam_depth*16+43)],data_in[`VWidth*(`APPRam_depth*15+44)-1:`VWidth*(`APPRam_depth*15+43)],data_in[`VWidth*(`APPRam_depth*14+44)-1:`VWidth*(`APPRam_depth*14+43)],data_in[`VWidth*(`APPRam_depth*13+44)-1:`VWidth*(`APPRam_depth*13+43)],data_in[`VWidth*(`APPRam_depth*12+44)-1:`VWidth*(`APPRam_depth*12+43)],data_in[`VWidth*(`APPRam_depth*11+44)-1:`VWidth*(`APPRam_depth*11+43)],data_in[`VWidth*(`APPRam_depth*10+44)-1:`VWidth*(`APPRam_depth*10+43)],data_in[`VWidth*(`APPRam_depth*9+44)-1:`VWidth*(`APPRam_depth*9+43)],data_in[`VWidth*(`APPRam_depth*8+44)-1:`VWidth*(`APPRam_depth*8+43)],data_in[`VWidth*(`APPRam_depth*7+44)-1:`VWidth*(`APPRam_depth*7+43)],data_in[`VWidth*(`APPRam_depth*6+44)-1:`VWidth*(`APPRam_depth*6+43)],data_in[`VWidth*(`APPRam_depth*5+44)-1:`VWidth*(`APPRam_depth*5+43)],data_in[`VWidth*(`APPRam_depth*4+44)-1:`VWidth*(`APPRam_depth*4+43)],data_in[`VWidth*(`APPRam_depth*3+44)-1:`VWidth*(`APPRam_depth*3+43)],data_in[`VWidth*(`APPRam_depth*2+44)-1:`VWidth*(`APPRam_depth*2+43)],data_in[`VWidth*(`APPRam_depth*1+44)-1:`VWidth*(`APPRam_depth*1+43)],data_in[`VWidth*(`APPRam_depth*0+44)-1:`VWidth*(`APPRam_depth*0+43)]};
			end
			44:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+45)-1:`VWidth*(`APPRam_depth*31+44)],data_in[`VWidth*(`APPRam_depth*30+45)-1:`VWidth*(`APPRam_depth*30+44)],data_in[`VWidth*(`APPRam_depth*29+45)-1:`VWidth*(`APPRam_depth*29+44)],data_in[`VWidth*(`APPRam_depth*28+45)-1:`VWidth*(`APPRam_depth*28+44)],data_in[`VWidth*(`APPRam_depth*27+45)-1:`VWidth*(`APPRam_depth*27+44)],data_in[`VWidth*(`APPRam_depth*26+45)-1:`VWidth*(`APPRam_depth*26+44)],data_in[`VWidth*(`APPRam_depth*25+45)-1:`VWidth*(`APPRam_depth*25+44)],data_in[`VWidth*(`APPRam_depth*24+45)-1:`VWidth*(`APPRam_depth*24+44)],data_in[`VWidth*(`APPRam_depth*23+45)-1:`VWidth*(`APPRam_depth*23+44)],data_in[`VWidth*(`APPRam_depth*22+45)-1:`VWidth*(`APPRam_depth*22+44)],data_in[`VWidth*(`APPRam_depth*21+45)-1:`VWidth*(`APPRam_depth*21+44)],data_in[`VWidth*(`APPRam_depth*20+45)-1:`VWidth*(`APPRam_depth*20+44)],data_in[`VWidth*(`APPRam_depth*19+45)-1:`VWidth*(`APPRam_depth*19+44)],data_in[`VWidth*(`APPRam_depth*18+45)-1:`VWidth*(`APPRam_depth*18+44)],data_in[`VWidth*(`APPRam_depth*17+45)-1:`VWidth*(`APPRam_depth*17+44)],data_in[`VWidth*(`APPRam_depth*16+45)-1:`VWidth*(`APPRam_depth*16+44)],data_in[`VWidth*(`APPRam_depth*15+45)-1:`VWidth*(`APPRam_depth*15+44)],data_in[`VWidth*(`APPRam_depth*14+45)-1:`VWidth*(`APPRam_depth*14+44)],data_in[`VWidth*(`APPRam_depth*13+45)-1:`VWidth*(`APPRam_depth*13+44)],data_in[`VWidth*(`APPRam_depth*12+45)-1:`VWidth*(`APPRam_depth*12+44)],data_in[`VWidth*(`APPRam_depth*11+45)-1:`VWidth*(`APPRam_depth*11+44)],data_in[`VWidth*(`APPRam_depth*10+45)-1:`VWidth*(`APPRam_depth*10+44)],data_in[`VWidth*(`APPRam_depth*9+45)-1:`VWidth*(`APPRam_depth*9+44)],data_in[`VWidth*(`APPRam_depth*8+45)-1:`VWidth*(`APPRam_depth*8+44)],data_in[`VWidth*(`APPRam_depth*7+45)-1:`VWidth*(`APPRam_depth*7+44)],data_in[`VWidth*(`APPRam_depth*6+45)-1:`VWidth*(`APPRam_depth*6+44)],data_in[`VWidth*(`APPRam_depth*5+45)-1:`VWidth*(`APPRam_depth*5+44)],data_in[`VWidth*(`APPRam_depth*4+45)-1:`VWidth*(`APPRam_depth*4+44)],data_in[`VWidth*(`APPRam_depth*3+45)-1:`VWidth*(`APPRam_depth*3+44)],data_in[`VWidth*(`APPRam_depth*2+45)-1:`VWidth*(`APPRam_depth*2+44)],data_in[`VWidth*(`APPRam_depth*1+45)-1:`VWidth*(`APPRam_depth*1+44)],data_in[`VWidth*(`APPRam_depth*0+45)-1:`VWidth*(`APPRam_depth*0+44)]};
			end
			45:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+46)-1:`VWidth*(`APPRam_depth*31+45)],data_in[`VWidth*(`APPRam_depth*30+46)-1:`VWidth*(`APPRam_depth*30+45)],data_in[`VWidth*(`APPRam_depth*29+46)-1:`VWidth*(`APPRam_depth*29+45)],data_in[`VWidth*(`APPRam_depth*28+46)-1:`VWidth*(`APPRam_depth*28+45)],data_in[`VWidth*(`APPRam_depth*27+46)-1:`VWidth*(`APPRam_depth*27+45)],data_in[`VWidth*(`APPRam_depth*26+46)-1:`VWidth*(`APPRam_depth*26+45)],data_in[`VWidth*(`APPRam_depth*25+46)-1:`VWidth*(`APPRam_depth*25+45)],data_in[`VWidth*(`APPRam_depth*24+46)-1:`VWidth*(`APPRam_depth*24+45)],data_in[`VWidth*(`APPRam_depth*23+46)-1:`VWidth*(`APPRam_depth*23+45)],data_in[`VWidth*(`APPRam_depth*22+46)-1:`VWidth*(`APPRam_depth*22+45)],data_in[`VWidth*(`APPRam_depth*21+46)-1:`VWidth*(`APPRam_depth*21+45)],data_in[`VWidth*(`APPRam_depth*20+46)-1:`VWidth*(`APPRam_depth*20+45)],data_in[`VWidth*(`APPRam_depth*19+46)-1:`VWidth*(`APPRam_depth*19+45)],data_in[`VWidth*(`APPRam_depth*18+46)-1:`VWidth*(`APPRam_depth*18+45)],data_in[`VWidth*(`APPRam_depth*17+46)-1:`VWidth*(`APPRam_depth*17+45)],data_in[`VWidth*(`APPRam_depth*16+46)-1:`VWidth*(`APPRam_depth*16+45)],data_in[`VWidth*(`APPRam_depth*15+46)-1:`VWidth*(`APPRam_depth*15+45)],data_in[`VWidth*(`APPRam_depth*14+46)-1:`VWidth*(`APPRam_depth*14+45)],data_in[`VWidth*(`APPRam_depth*13+46)-1:`VWidth*(`APPRam_depth*13+45)],data_in[`VWidth*(`APPRam_depth*12+46)-1:`VWidth*(`APPRam_depth*12+45)],data_in[`VWidth*(`APPRam_depth*11+46)-1:`VWidth*(`APPRam_depth*11+45)],data_in[`VWidth*(`APPRam_depth*10+46)-1:`VWidth*(`APPRam_depth*10+45)],data_in[`VWidth*(`APPRam_depth*9+46)-1:`VWidth*(`APPRam_depth*9+45)],data_in[`VWidth*(`APPRam_depth*8+46)-1:`VWidth*(`APPRam_depth*8+45)],data_in[`VWidth*(`APPRam_depth*7+46)-1:`VWidth*(`APPRam_depth*7+45)],data_in[`VWidth*(`APPRam_depth*6+46)-1:`VWidth*(`APPRam_depth*6+45)],data_in[`VWidth*(`APPRam_depth*5+46)-1:`VWidth*(`APPRam_depth*5+45)],data_in[`VWidth*(`APPRam_depth*4+46)-1:`VWidth*(`APPRam_depth*4+45)],data_in[`VWidth*(`APPRam_depth*3+46)-1:`VWidth*(`APPRam_depth*3+45)],data_in[`VWidth*(`APPRam_depth*2+46)-1:`VWidth*(`APPRam_depth*2+45)],data_in[`VWidth*(`APPRam_depth*1+46)-1:`VWidth*(`APPRam_depth*1+45)],data_in[`VWidth*(`APPRam_depth*0+46)-1:`VWidth*(`APPRam_depth*0+45)]};
			end
			46:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+47)-1:`VWidth*(`APPRam_depth*31+46)],data_in[`VWidth*(`APPRam_depth*30+47)-1:`VWidth*(`APPRam_depth*30+46)],data_in[`VWidth*(`APPRam_depth*29+47)-1:`VWidth*(`APPRam_depth*29+46)],data_in[`VWidth*(`APPRam_depth*28+47)-1:`VWidth*(`APPRam_depth*28+46)],data_in[`VWidth*(`APPRam_depth*27+47)-1:`VWidth*(`APPRam_depth*27+46)],data_in[`VWidth*(`APPRam_depth*26+47)-1:`VWidth*(`APPRam_depth*26+46)],data_in[`VWidth*(`APPRam_depth*25+47)-1:`VWidth*(`APPRam_depth*25+46)],data_in[`VWidth*(`APPRam_depth*24+47)-1:`VWidth*(`APPRam_depth*24+46)],data_in[`VWidth*(`APPRam_depth*23+47)-1:`VWidth*(`APPRam_depth*23+46)],data_in[`VWidth*(`APPRam_depth*22+47)-1:`VWidth*(`APPRam_depth*22+46)],data_in[`VWidth*(`APPRam_depth*21+47)-1:`VWidth*(`APPRam_depth*21+46)],data_in[`VWidth*(`APPRam_depth*20+47)-1:`VWidth*(`APPRam_depth*20+46)],data_in[`VWidth*(`APPRam_depth*19+47)-1:`VWidth*(`APPRam_depth*19+46)],data_in[`VWidth*(`APPRam_depth*18+47)-1:`VWidth*(`APPRam_depth*18+46)],data_in[`VWidth*(`APPRam_depth*17+47)-1:`VWidth*(`APPRam_depth*17+46)],data_in[`VWidth*(`APPRam_depth*16+47)-1:`VWidth*(`APPRam_depth*16+46)],data_in[`VWidth*(`APPRam_depth*15+47)-1:`VWidth*(`APPRam_depth*15+46)],data_in[`VWidth*(`APPRam_depth*14+47)-1:`VWidth*(`APPRam_depth*14+46)],data_in[`VWidth*(`APPRam_depth*13+47)-1:`VWidth*(`APPRam_depth*13+46)],data_in[`VWidth*(`APPRam_depth*12+47)-1:`VWidth*(`APPRam_depth*12+46)],data_in[`VWidth*(`APPRam_depth*11+47)-1:`VWidth*(`APPRam_depth*11+46)],data_in[`VWidth*(`APPRam_depth*10+47)-1:`VWidth*(`APPRam_depth*10+46)],data_in[`VWidth*(`APPRam_depth*9+47)-1:`VWidth*(`APPRam_depth*9+46)],data_in[`VWidth*(`APPRam_depth*8+47)-1:`VWidth*(`APPRam_depth*8+46)],data_in[`VWidth*(`APPRam_depth*7+47)-1:`VWidth*(`APPRam_depth*7+46)],data_in[`VWidth*(`APPRam_depth*6+47)-1:`VWidth*(`APPRam_depth*6+46)],data_in[`VWidth*(`APPRam_depth*5+47)-1:`VWidth*(`APPRam_depth*5+46)],data_in[`VWidth*(`APPRam_depth*4+47)-1:`VWidth*(`APPRam_depth*4+46)],data_in[`VWidth*(`APPRam_depth*3+47)-1:`VWidth*(`APPRam_depth*3+46)],data_in[`VWidth*(`APPRam_depth*2+47)-1:`VWidth*(`APPRam_depth*2+46)],data_in[`VWidth*(`APPRam_depth*1+47)-1:`VWidth*(`APPRam_depth*1+46)],data_in[`VWidth*(`APPRam_depth*0+47)-1:`VWidth*(`APPRam_depth*0+46)]};
			end
			47:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+48)-1:`VWidth*(`APPRam_depth*31+47)],data_in[`VWidth*(`APPRam_depth*30+48)-1:`VWidth*(`APPRam_depth*30+47)],data_in[`VWidth*(`APPRam_depth*29+48)-1:`VWidth*(`APPRam_depth*29+47)],data_in[`VWidth*(`APPRam_depth*28+48)-1:`VWidth*(`APPRam_depth*28+47)],data_in[`VWidth*(`APPRam_depth*27+48)-1:`VWidth*(`APPRam_depth*27+47)],data_in[`VWidth*(`APPRam_depth*26+48)-1:`VWidth*(`APPRam_depth*26+47)],data_in[`VWidth*(`APPRam_depth*25+48)-1:`VWidth*(`APPRam_depth*25+47)],data_in[`VWidth*(`APPRam_depth*24+48)-1:`VWidth*(`APPRam_depth*24+47)],data_in[`VWidth*(`APPRam_depth*23+48)-1:`VWidth*(`APPRam_depth*23+47)],data_in[`VWidth*(`APPRam_depth*22+48)-1:`VWidth*(`APPRam_depth*22+47)],data_in[`VWidth*(`APPRam_depth*21+48)-1:`VWidth*(`APPRam_depth*21+47)],data_in[`VWidth*(`APPRam_depth*20+48)-1:`VWidth*(`APPRam_depth*20+47)],data_in[`VWidth*(`APPRam_depth*19+48)-1:`VWidth*(`APPRam_depth*19+47)],data_in[`VWidth*(`APPRam_depth*18+48)-1:`VWidth*(`APPRam_depth*18+47)],data_in[`VWidth*(`APPRam_depth*17+48)-1:`VWidth*(`APPRam_depth*17+47)],data_in[`VWidth*(`APPRam_depth*16+48)-1:`VWidth*(`APPRam_depth*16+47)],data_in[`VWidth*(`APPRam_depth*15+48)-1:`VWidth*(`APPRam_depth*15+47)],data_in[`VWidth*(`APPRam_depth*14+48)-1:`VWidth*(`APPRam_depth*14+47)],data_in[`VWidth*(`APPRam_depth*13+48)-1:`VWidth*(`APPRam_depth*13+47)],data_in[`VWidth*(`APPRam_depth*12+48)-1:`VWidth*(`APPRam_depth*12+47)],data_in[`VWidth*(`APPRam_depth*11+48)-1:`VWidth*(`APPRam_depth*11+47)],data_in[`VWidth*(`APPRam_depth*10+48)-1:`VWidth*(`APPRam_depth*10+47)],data_in[`VWidth*(`APPRam_depth*9+48)-1:`VWidth*(`APPRam_depth*9+47)],data_in[`VWidth*(`APPRam_depth*8+48)-1:`VWidth*(`APPRam_depth*8+47)],data_in[`VWidth*(`APPRam_depth*7+48)-1:`VWidth*(`APPRam_depth*7+47)],data_in[`VWidth*(`APPRam_depth*6+48)-1:`VWidth*(`APPRam_depth*6+47)],data_in[`VWidth*(`APPRam_depth*5+48)-1:`VWidth*(`APPRam_depth*5+47)],data_in[`VWidth*(`APPRam_depth*4+48)-1:`VWidth*(`APPRam_depth*4+47)],data_in[`VWidth*(`APPRam_depth*3+48)-1:`VWidth*(`APPRam_depth*3+47)],data_in[`VWidth*(`APPRam_depth*2+48)-1:`VWidth*(`APPRam_depth*2+47)],data_in[`VWidth*(`APPRam_depth*1+48)-1:`VWidth*(`APPRam_depth*1+47)],data_in[`VWidth*(`APPRam_depth*0+48)-1:`VWidth*(`APPRam_depth*0+47)]};
			end
			48:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+49)-1:`VWidth*(`APPRam_depth*31+48)],data_in[`VWidth*(`APPRam_depth*30+49)-1:`VWidth*(`APPRam_depth*30+48)],data_in[`VWidth*(`APPRam_depth*29+49)-1:`VWidth*(`APPRam_depth*29+48)],data_in[`VWidth*(`APPRam_depth*28+49)-1:`VWidth*(`APPRam_depth*28+48)],data_in[`VWidth*(`APPRam_depth*27+49)-1:`VWidth*(`APPRam_depth*27+48)],data_in[`VWidth*(`APPRam_depth*26+49)-1:`VWidth*(`APPRam_depth*26+48)],data_in[`VWidth*(`APPRam_depth*25+49)-1:`VWidth*(`APPRam_depth*25+48)],data_in[`VWidth*(`APPRam_depth*24+49)-1:`VWidth*(`APPRam_depth*24+48)],data_in[`VWidth*(`APPRam_depth*23+49)-1:`VWidth*(`APPRam_depth*23+48)],data_in[`VWidth*(`APPRam_depth*22+49)-1:`VWidth*(`APPRam_depth*22+48)],data_in[`VWidth*(`APPRam_depth*21+49)-1:`VWidth*(`APPRam_depth*21+48)],data_in[`VWidth*(`APPRam_depth*20+49)-1:`VWidth*(`APPRam_depth*20+48)],data_in[`VWidth*(`APPRam_depth*19+49)-1:`VWidth*(`APPRam_depth*19+48)],data_in[`VWidth*(`APPRam_depth*18+49)-1:`VWidth*(`APPRam_depth*18+48)],data_in[`VWidth*(`APPRam_depth*17+49)-1:`VWidth*(`APPRam_depth*17+48)],data_in[`VWidth*(`APPRam_depth*16+49)-1:`VWidth*(`APPRam_depth*16+48)],data_in[`VWidth*(`APPRam_depth*15+49)-1:`VWidth*(`APPRam_depth*15+48)],data_in[`VWidth*(`APPRam_depth*14+49)-1:`VWidth*(`APPRam_depth*14+48)],data_in[`VWidth*(`APPRam_depth*13+49)-1:`VWidth*(`APPRam_depth*13+48)],data_in[`VWidth*(`APPRam_depth*12+49)-1:`VWidth*(`APPRam_depth*12+48)],data_in[`VWidth*(`APPRam_depth*11+49)-1:`VWidth*(`APPRam_depth*11+48)],data_in[`VWidth*(`APPRam_depth*10+49)-1:`VWidth*(`APPRam_depth*10+48)],data_in[`VWidth*(`APPRam_depth*9+49)-1:`VWidth*(`APPRam_depth*9+48)],data_in[`VWidth*(`APPRam_depth*8+49)-1:`VWidth*(`APPRam_depth*8+48)],data_in[`VWidth*(`APPRam_depth*7+49)-1:`VWidth*(`APPRam_depth*7+48)],data_in[`VWidth*(`APPRam_depth*6+49)-1:`VWidth*(`APPRam_depth*6+48)],data_in[`VWidth*(`APPRam_depth*5+49)-1:`VWidth*(`APPRam_depth*5+48)],data_in[`VWidth*(`APPRam_depth*4+49)-1:`VWidth*(`APPRam_depth*4+48)],data_in[`VWidth*(`APPRam_depth*3+49)-1:`VWidth*(`APPRam_depth*3+48)],data_in[`VWidth*(`APPRam_depth*2+49)-1:`VWidth*(`APPRam_depth*2+48)],data_in[`VWidth*(`APPRam_depth*1+49)-1:`VWidth*(`APPRam_depth*1+48)],data_in[`VWidth*(`APPRam_depth*0+49)-1:`VWidth*(`APPRam_depth*0+48)]};
			end
			49:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+50)-1:`VWidth*(`APPRam_depth*31+49)],data_in[`VWidth*(`APPRam_depth*30+50)-1:`VWidth*(`APPRam_depth*30+49)],data_in[`VWidth*(`APPRam_depth*29+50)-1:`VWidth*(`APPRam_depth*29+49)],data_in[`VWidth*(`APPRam_depth*28+50)-1:`VWidth*(`APPRam_depth*28+49)],data_in[`VWidth*(`APPRam_depth*27+50)-1:`VWidth*(`APPRam_depth*27+49)],data_in[`VWidth*(`APPRam_depth*26+50)-1:`VWidth*(`APPRam_depth*26+49)],data_in[`VWidth*(`APPRam_depth*25+50)-1:`VWidth*(`APPRam_depth*25+49)],data_in[`VWidth*(`APPRam_depth*24+50)-1:`VWidth*(`APPRam_depth*24+49)],data_in[`VWidth*(`APPRam_depth*23+50)-1:`VWidth*(`APPRam_depth*23+49)],data_in[`VWidth*(`APPRam_depth*22+50)-1:`VWidth*(`APPRam_depth*22+49)],data_in[`VWidth*(`APPRam_depth*21+50)-1:`VWidth*(`APPRam_depth*21+49)],data_in[`VWidth*(`APPRam_depth*20+50)-1:`VWidth*(`APPRam_depth*20+49)],data_in[`VWidth*(`APPRam_depth*19+50)-1:`VWidth*(`APPRam_depth*19+49)],data_in[`VWidth*(`APPRam_depth*18+50)-1:`VWidth*(`APPRam_depth*18+49)],data_in[`VWidth*(`APPRam_depth*17+50)-1:`VWidth*(`APPRam_depth*17+49)],data_in[`VWidth*(`APPRam_depth*16+50)-1:`VWidth*(`APPRam_depth*16+49)],data_in[`VWidth*(`APPRam_depth*15+50)-1:`VWidth*(`APPRam_depth*15+49)],data_in[`VWidth*(`APPRam_depth*14+50)-1:`VWidth*(`APPRam_depth*14+49)],data_in[`VWidth*(`APPRam_depth*13+50)-1:`VWidth*(`APPRam_depth*13+49)],data_in[`VWidth*(`APPRam_depth*12+50)-1:`VWidth*(`APPRam_depth*12+49)],data_in[`VWidth*(`APPRam_depth*11+50)-1:`VWidth*(`APPRam_depth*11+49)],data_in[`VWidth*(`APPRam_depth*10+50)-1:`VWidth*(`APPRam_depth*10+49)],data_in[`VWidth*(`APPRam_depth*9+50)-1:`VWidth*(`APPRam_depth*9+49)],data_in[`VWidth*(`APPRam_depth*8+50)-1:`VWidth*(`APPRam_depth*8+49)],data_in[`VWidth*(`APPRam_depth*7+50)-1:`VWidth*(`APPRam_depth*7+49)],data_in[`VWidth*(`APPRam_depth*6+50)-1:`VWidth*(`APPRam_depth*6+49)],data_in[`VWidth*(`APPRam_depth*5+50)-1:`VWidth*(`APPRam_depth*5+49)],data_in[`VWidth*(`APPRam_depth*4+50)-1:`VWidth*(`APPRam_depth*4+49)],data_in[`VWidth*(`APPRam_depth*3+50)-1:`VWidth*(`APPRam_depth*3+49)],data_in[`VWidth*(`APPRam_depth*2+50)-1:`VWidth*(`APPRam_depth*2+49)],data_in[`VWidth*(`APPRam_depth*1+50)-1:`VWidth*(`APPRam_depth*1+49)],data_in[`VWidth*(`APPRam_depth*0+50)-1:`VWidth*(`APPRam_depth*0+49)]};
			end
			50:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+51)-1:`VWidth*(`APPRam_depth*31+50)],data_in[`VWidth*(`APPRam_depth*30+51)-1:`VWidth*(`APPRam_depth*30+50)],data_in[`VWidth*(`APPRam_depth*29+51)-1:`VWidth*(`APPRam_depth*29+50)],data_in[`VWidth*(`APPRam_depth*28+51)-1:`VWidth*(`APPRam_depth*28+50)],data_in[`VWidth*(`APPRam_depth*27+51)-1:`VWidth*(`APPRam_depth*27+50)],data_in[`VWidth*(`APPRam_depth*26+51)-1:`VWidth*(`APPRam_depth*26+50)],data_in[`VWidth*(`APPRam_depth*25+51)-1:`VWidth*(`APPRam_depth*25+50)],data_in[`VWidth*(`APPRam_depth*24+51)-1:`VWidth*(`APPRam_depth*24+50)],data_in[`VWidth*(`APPRam_depth*23+51)-1:`VWidth*(`APPRam_depth*23+50)],data_in[`VWidth*(`APPRam_depth*22+51)-1:`VWidth*(`APPRam_depth*22+50)],data_in[`VWidth*(`APPRam_depth*21+51)-1:`VWidth*(`APPRam_depth*21+50)],data_in[`VWidth*(`APPRam_depth*20+51)-1:`VWidth*(`APPRam_depth*20+50)],data_in[`VWidth*(`APPRam_depth*19+51)-1:`VWidth*(`APPRam_depth*19+50)],data_in[`VWidth*(`APPRam_depth*18+51)-1:`VWidth*(`APPRam_depth*18+50)],data_in[`VWidth*(`APPRam_depth*17+51)-1:`VWidth*(`APPRam_depth*17+50)],data_in[`VWidth*(`APPRam_depth*16+51)-1:`VWidth*(`APPRam_depth*16+50)],data_in[`VWidth*(`APPRam_depth*15+51)-1:`VWidth*(`APPRam_depth*15+50)],data_in[`VWidth*(`APPRam_depth*14+51)-1:`VWidth*(`APPRam_depth*14+50)],data_in[`VWidth*(`APPRam_depth*13+51)-1:`VWidth*(`APPRam_depth*13+50)],data_in[`VWidth*(`APPRam_depth*12+51)-1:`VWidth*(`APPRam_depth*12+50)],data_in[`VWidth*(`APPRam_depth*11+51)-1:`VWidth*(`APPRam_depth*11+50)],data_in[`VWidth*(`APPRam_depth*10+51)-1:`VWidth*(`APPRam_depth*10+50)],data_in[`VWidth*(`APPRam_depth*9+51)-1:`VWidth*(`APPRam_depth*9+50)],data_in[`VWidth*(`APPRam_depth*8+51)-1:`VWidth*(`APPRam_depth*8+50)],data_in[`VWidth*(`APPRam_depth*7+51)-1:`VWidth*(`APPRam_depth*7+50)],data_in[`VWidth*(`APPRam_depth*6+51)-1:`VWidth*(`APPRam_depth*6+50)],data_in[`VWidth*(`APPRam_depth*5+51)-1:`VWidth*(`APPRam_depth*5+50)],data_in[`VWidth*(`APPRam_depth*4+51)-1:`VWidth*(`APPRam_depth*4+50)],data_in[`VWidth*(`APPRam_depth*3+51)-1:`VWidth*(`APPRam_depth*3+50)],data_in[`VWidth*(`APPRam_depth*2+51)-1:`VWidth*(`APPRam_depth*2+50)],data_in[`VWidth*(`APPRam_depth*1+51)-1:`VWidth*(`APPRam_depth*1+50)],data_in[`VWidth*(`APPRam_depth*0+51)-1:`VWidth*(`APPRam_depth*0+50)]};
			end
			51:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+52)-1:`VWidth*(`APPRam_depth*31+51)],data_in[`VWidth*(`APPRam_depth*30+52)-1:`VWidth*(`APPRam_depth*30+51)],data_in[`VWidth*(`APPRam_depth*29+52)-1:`VWidth*(`APPRam_depth*29+51)],data_in[`VWidth*(`APPRam_depth*28+52)-1:`VWidth*(`APPRam_depth*28+51)],data_in[`VWidth*(`APPRam_depth*27+52)-1:`VWidth*(`APPRam_depth*27+51)],data_in[`VWidth*(`APPRam_depth*26+52)-1:`VWidth*(`APPRam_depth*26+51)],data_in[`VWidth*(`APPRam_depth*25+52)-1:`VWidth*(`APPRam_depth*25+51)],data_in[`VWidth*(`APPRam_depth*24+52)-1:`VWidth*(`APPRam_depth*24+51)],data_in[`VWidth*(`APPRam_depth*23+52)-1:`VWidth*(`APPRam_depth*23+51)],data_in[`VWidth*(`APPRam_depth*22+52)-1:`VWidth*(`APPRam_depth*22+51)],data_in[`VWidth*(`APPRam_depth*21+52)-1:`VWidth*(`APPRam_depth*21+51)],data_in[`VWidth*(`APPRam_depth*20+52)-1:`VWidth*(`APPRam_depth*20+51)],data_in[`VWidth*(`APPRam_depth*19+52)-1:`VWidth*(`APPRam_depth*19+51)],data_in[`VWidth*(`APPRam_depth*18+52)-1:`VWidth*(`APPRam_depth*18+51)],data_in[`VWidth*(`APPRam_depth*17+52)-1:`VWidth*(`APPRam_depth*17+51)],data_in[`VWidth*(`APPRam_depth*16+52)-1:`VWidth*(`APPRam_depth*16+51)],data_in[`VWidth*(`APPRam_depth*15+52)-1:`VWidth*(`APPRam_depth*15+51)],data_in[`VWidth*(`APPRam_depth*14+52)-1:`VWidth*(`APPRam_depth*14+51)],data_in[`VWidth*(`APPRam_depth*13+52)-1:`VWidth*(`APPRam_depth*13+51)],data_in[`VWidth*(`APPRam_depth*12+52)-1:`VWidth*(`APPRam_depth*12+51)],data_in[`VWidth*(`APPRam_depth*11+52)-1:`VWidth*(`APPRam_depth*11+51)],data_in[`VWidth*(`APPRam_depth*10+52)-1:`VWidth*(`APPRam_depth*10+51)],data_in[`VWidth*(`APPRam_depth*9+52)-1:`VWidth*(`APPRam_depth*9+51)],data_in[`VWidth*(`APPRam_depth*8+52)-1:`VWidth*(`APPRam_depth*8+51)],data_in[`VWidth*(`APPRam_depth*7+52)-1:`VWidth*(`APPRam_depth*7+51)],data_in[`VWidth*(`APPRam_depth*6+52)-1:`VWidth*(`APPRam_depth*6+51)],data_in[`VWidth*(`APPRam_depth*5+52)-1:`VWidth*(`APPRam_depth*5+51)],data_in[`VWidth*(`APPRam_depth*4+52)-1:`VWidth*(`APPRam_depth*4+51)],data_in[`VWidth*(`APPRam_depth*3+52)-1:`VWidth*(`APPRam_depth*3+51)],data_in[`VWidth*(`APPRam_depth*2+52)-1:`VWidth*(`APPRam_depth*2+51)],data_in[`VWidth*(`APPRam_depth*1+52)-1:`VWidth*(`APPRam_depth*1+51)],data_in[`VWidth*(`APPRam_depth*0+52)-1:`VWidth*(`APPRam_depth*0+51)]};
			end
			52:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+53)-1:`VWidth*(`APPRam_depth*31+52)],data_in[`VWidth*(`APPRam_depth*30+53)-1:`VWidth*(`APPRam_depth*30+52)],data_in[`VWidth*(`APPRam_depth*29+53)-1:`VWidth*(`APPRam_depth*29+52)],data_in[`VWidth*(`APPRam_depth*28+53)-1:`VWidth*(`APPRam_depth*28+52)],data_in[`VWidth*(`APPRam_depth*27+53)-1:`VWidth*(`APPRam_depth*27+52)],data_in[`VWidth*(`APPRam_depth*26+53)-1:`VWidth*(`APPRam_depth*26+52)],data_in[`VWidth*(`APPRam_depth*25+53)-1:`VWidth*(`APPRam_depth*25+52)],data_in[`VWidth*(`APPRam_depth*24+53)-1:`VWidth*(`APPRam_depth*24+52)],data_in[`VWidth*(`APPRam_depth*23+53)-1:`VWidth*(`APPRam_depth*23+52)],data_in[`VWidth*(`APPRam_depth*22+53)-1:`VWidth*(`APPRam_depth*22+52)],data_in[`VWidth*(`APPRam_depth*21+53)-1:`VWidth*(`APPRam_depth*21+52)],data_in[`VWidth*(`APPRam_depth*20+53)-1:`VWidth*(`APPRam_depth*20+52)],data_in[`VWidth*(`APPRam_depth*19+53)-1:`VWidth*(`APPRam_depth*19+52)],data_in[`VWidth*(`APPRam_depth*18+53)-1:`VWidth*(`APPRam_depth*18+52)],data_in[`VWidth*(`APPRam_depth*17+53)-1:`VWidth*(`APPRam_depth*17+52)],data_in[`VWidth*(`APPRam_depth*16+53)-1:`VWidth*(`APPRam_depth*16+52)],data_in[`VWidth*(`APPRam_depth*15+53)-1:`VWidth*(`APPRam_depth*15+52)],data_in[`VWidth*(`APPRam_depth*14+53)-1:`VWidth*(`APPRam_depth*14+52)],data_in[`VWidth*(`APPRam_depth*13+53)-1:`VWidth*(`APPRam_depth*13+52)],data_in[`VWidth*(`APPRam_depth*12+53)-1:`VWidth*(`APPRam_depth*12+52)],data_in[`VWidth*(`APPRam_depth*11+53)-1:`VWidth*(`APPRam_depth*11+52)],data_in[`VWidth*(`APPRam_depth*10+53)-1:`VWidth*(`APPRam_depth*10+52)],data_in[`VWidth*(`APPRam_depth*9+53)-1:`VWidth*(`APPRam_depth*9+52)],data_in[`VWidth*(`APPRam_depth*8+53)-1:`VWidth*(`APPRam_depth*8+52)],data_in[`VWidth*(`APPRam_depth*7+53)-1:`VWidth*(`APPRam_depth*7+52)],data_in[`VWidth*(`APPRam_depth*6+53)-1:`VWidth*(`APPRam_depth*6+52)],data_in[`VWidth*(`APPRam_depth*5+53)-1:`VWidth*(`APPRam_depth*5+52)],data_in[`VWidth*(`APPRam_depth*4+53)-1:`VWidth*(`APPRam_depth*4+52)],data_in[`VWidth*(`APPRam_depth*3+53)-1:`VWidth*(`APPRam_depth*3+52)],data_in[`VWidth*(`APPRam_depth*2+53)-1:`VWidth*(`APPRam_depth*2+52)],data_in[`VWidth*(`APPRam_depth*1+53)-1:`VWidth*(`APPRam_depth*1+52)],data_in[`VWidth*(`APPRam_depth*0+53)-1:`VWidth*(`APPRam_depth*0+52)]};
			end
			53:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+54)-1:`VWidth*(`APPRam_depth*31+53)],data_in[`VWidth*(`APPRam_depth*30+54)-1:`VWidth*(`APPRam_depth*30+53)],data_in[`VWidth*(`APPRam_depth*29+54)-1:`VWidth*(`APPRam_depth*29+53)],data_in[`VWidth*(`APPRam_depth*28+54)-1:`VWidth*(`APPRam_depth*28+53)],data_in[`VWidth*(`APPRam_depth*27+54)-1:`VWidth*(`APPRam_depth*27+53)],data_in[`VWidth*(`APPRam_depth*26+54)-1:`VWidth*(`APPRam_depth*26+53)],data_in[`VWidth*(`APPRam_depth*25+54)-1:`VWidth*(`APPRam_depth*25+53)],data_in[`VWidth*(`APPRam_depth*24+54)-1:`VWidth*(`APPRam_depth*24+53)],data_in[`VWidth*(`APPRam_depth*23+54)-1:`VWidth*(`APPRam_depth*23+53)],data_in[`VWidth*(`APPRam_depth*22+54)-1:`VWidth*(`APPRam_depth*22+53)],data_in[`VWidth*(`APPRam_depth*21+54)-1:`VWidth*(`APPRam_depth*21+53)],data_in[`VWidth*(`APPRam_depth*20+54)-1:`VWidth*(`APPRam_depth*20+53)],data_in[`VWidth*(`APPRam_depth*19+54)-1:`VWidth*(`APPRam_depth*19+53)],data_in[`VWidth*(`APPRam_depth*18+54)-1:`VWidth*(`APPRam_depth*18+53)],data_in[`VWidth*(`APPRam_depth*17+54)-1:`VWidth*(`APPRam_depth*17+53)],data_in[`VWidth*(`APPRam_depth*16+54)-1:`VWidth*(`APPRam_depth*16+53)],data_in[`VWidth*(`APPRam_depth*15+54)-1:`VWidth*(`APPRam_depth*15+53)],data_in[`VWidth*(`APPRam_depth*14+54)-1:`VWidth*(`APPRam_depth*14+53)],data_in[`VWidth*(`APPRam_depth*13+54)-1:`VWidth*(`APPRam_depth*13+53)],data_in[`VWidth*(`APPRam_depth*12+54)-1:`VWidth*(`APPRam_depth*12+53)],data_in[`VWidth*(`APPRam_depth*11+54)-1:`VWidth*(`APPRam_depth*11+53)],data_in[`VWidth*(`APPRam_depth*10+54)-1:`VWidth*(`APPRam_depth*10+53)],data_in[`VWidth*(`APPRam_depth*9+54)-1:`VWidth*(`APPRam_depth*9+53)],data_in[`VWidth*(`APPRam_depth*8+54)-1:`VWidth*(`APPRam_depth*8+53)],data_in[`VWidth*(`APPRam_depth*7+54)-1:`VWidth*(`APPRam_depth*7+53)],data_in[`VWidth*(`APPRam_depth*6+54)-1:`VWidth*(`APPRam_depth*6+53)],data_in[`VWidth*(`APPRam_depth*5+54)-1:`VWidth*(`APPRam_depth*5+53)],data_in[`VWidth*(`APPRam_depth*4+54)-1:`VWidth*(`APPRam_depth*4+53)],data_in[`VWidth*(`APPRam_depth*3+54)-1:`VWidth*(`APPRam_depth*3+53)],data_in[`VWidth*(`APPRam_depth*2+54)-1:`VWidth*(`APPRam_depth*2+53)],data_in[`VWidth*(`APPRam_depth*1+54)-1:`VWidth*(`APPRam_depth*1+53)],data_in[`VWidth*(`APPRam_depth*0+54)-1:`VWidth*(`APPRam_depth*0+53)]};
			end
			54:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+55)-1:`VWidth*(`APPRam_depth*31+54)],data_in[`VWidth*(`APPRam_depth*30+55)-1:`VWidth*(`APPRam_depth*30+54)],data_in[`VWidth*(`APPRam_depth*29+55)-1:`VWidth*(`APPRam_depth*29+54)],data_in[`VWidth*(`APPRam_depth*28+55)-1:`VWidth*(`APPRam_depth*28+54)],data_in[`VWidth*(`APPRam_depth*27+55)-1:`VWidth*(`APPRam_depth*27+54)],data_in[`VWidth*(`APPRam_depth*26+55)-1:`VWidth*(`APPRam_depth*26+54)],data_in[`VWidth*(`APPRam_depth*25+55)-1:`VWidth*(`APPRam_depth*25+54)],data_in[`VWidth*(`APPRam_depth*24+55)-1:`VWidth*(`APPRam_depth*24+54)],data_in[`VWidth*(`APPRam_depth*23+55)-1:`VWidth*(`APPRam_depth*23+54)],data_in[`VWidth*(`APPRam_depth*22+55)-1:`VWidth*(`APPRam_depth*22+54)],data_in[`VWidth*(`APPRam_depth*21+55)-1:`VWidth*(`APPRam_depth*21+54)],data_in[`VWidth*(`APPRam_depth*20+55)-1:`VWidth*(`APPRam_depth*20+54)],data_in[`VWidth*(`APPRam_depth*19+55)-1:`VWidth*(`APPRam_depth*19+54)],data_in[`VWidth*(`APPRam_depth*18+55)-1:`VWidth*(`APPRam_depth*18+54)],data_in[`VWidth*(`APPRam_depth*17+55)-1:`VWidth*(`APPRam_depth*17+54)],data_in[`VWidth*(`APPRam_depth*16+55)-1:`VWidth*(`APPRam_depth*16+54)],data_in[`VWidth*(`APPRam_depth*15+55)-1:`VWidth*(`APPRam_depth*15+54)],data_in[`VWidth*(`APPRam_depth*14+55)-1:`VWidth*(`APPRam_depth*14+54)],data_in[`VWidth*(`APPRam_depth*13+55)-1:`VWidth*(`APPRam_depth*13+54)],data_in[`VWidth*(`APPRam_depth*12+55)-1:`VWidth*(`APPRam_depth*12+54)],data_in[`VWidth*(`APPRam_depth*11+55)-1:`VWidth*(`APPRam_depth*11+54)],data_in[`VWidth*(`APPRam_depth*10+55)-1:`VWidth*(`APPRam_depth*10+54)],data_in[`VWidth*(`APPRam_depth*9+55)-1:`VWidth*(`APPRam_depth*9+54)],data_in[`VWidth*(`APPRam_depth*8+55)-1:`VWidth*(`APPRam_depth*8+54)],data_in[`VWidth*(`APPRam_depth*7+55)-1:`VWidth*(`APPRam_depth*7+54)],data_in[`VWidth*(`APPRam_depth*6+55)-1:`VWidth*(`APPRam_depth*6+54)],data_in[`VWidth*(`APPRam_depth*5+55)-1:`VWidth*(`APPRam_depth*5+54)],data_in[`VWidth*(`APPRam_depth*4+55)-1:`VWidth*(`APPRam_depth*4+54)],data_in[`VWidth*(`APPRam_depth*3+55)-1:`VWidth*(`APPRam_depth*3+54)],data_in[`VWidth*(`APPRam_depth*2+55)-1:`VWidth*(`APPRam_depth*2+54)],data_in[`VWidth*(`APPRam_depth*1+55)-1:`VWidth*(`APPRam_depth*1+54)],data_in[`VWidth*(`APPRam_depth*0+55)-1:`VWidth*(`APPRam_depth*0+54)]};
			end
			55:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+56)-1:`VWidth*(`APPRam_depth*31+55)],data_in[`VWidth*(`APPRam_depth*30+56)-1:`VWidth*(`APPRam_depth*30+55)],data_in[`VWidth*(`APPRam_depth*29+56)-1:`VWidth*(`APPRam_depth*29+55)],data_in[`VWidth*(`APPRam_depth*28+56)-1:`VWidth*(`APPRam_depth*28+55)],data_in[`VWidth*(`APPRam_depth*27+56)-1:`VWidth*(`APPRam_depth*27+55)],data_in[`VWidth*(`APPRam_depth*26+56)-1:`VWidth*(`APPRam_depth*26+55)],data_in[`VWidth*(`APPRam_depth*25+56)-1:`VWidth*(`APPRam_depth*25+55)],data_in[`VWidth*(`APPRam_depth*24+56)-1:`VWidth*(`APPRam_depth*24+55)],data_in[`VWidth*(`APPRam_depth*23+56)-1:`VWidth*(`APPRam_depth*23+55)],data_in[`VWidth*(`APPRam_depth*22+56)-1:`VWidth*(`APPRam_depth*22+55)],data_in[`VWidth*(`APPRam_depth*21+56)-1:`VWidth*(`APPRam_depth*21+55)],data_in[`VWidth*(`APPRam_depth*20+56)-1:`VWidth*(`APPRam_depth*20+55)],data_in[`VWidth*(`APPRam_depth*19+56)-1:`VWidth*(`APPRam_depth*19+55)],data_in[`VWidth*(`APPRam_depth*18+56)-1:`VWidth*(`APPRam_depth*18+55)],data_in[`VWidth*(`APPRam_depth*17+56)-1:`VWidth*(`APPRam_depth*17+55)],data_in[`VWidth*(`APPRam_depth*16+56)-1:`VWidth*(`APPRam_depth*16+55)],data_in[`VWidth*(`APPRam_depth*15+56)-1:`VWidth*(`APPRam_depth*15+55)],data_in[`VWidth*(`APPRam_depth*14+56)-1:`VWidth*(`APPRam_depth*14+55)],data_in[`VWidth*(`APPRam_depth*13+56)-1:`VWidth*(`APPRam_depth*13+55)],data_in[`VWidth*(`APPRam_depth*12+56)-1:`VWidth*(`APPRam_depth*12+55)],data_in[`VWidth*(`APPRam_depth*11+56)-1:`VWidth*(`APPRam_depth*11+55)],data_in[`VWidth*(`APPRam_depth*10+56)-1:`VWidth*(`APPRam_depth*10+55)],data_in[`VWidth*(`APPRam_depth*9+56)-1:`VWidth*(`APPRam_depth*9+55)],data_in[`VWidth*(`APPRam_depth*8+56)-1:`VWidth*(`APPRam_depth*8+55)],data_in[`VWidth*(`APPRam_depth*7+56)-1:`VWidth*(`APPRam_depth*7+55)],data_in[`VWidth*(`APPRam_depth*6+56)-1:`VWidth*(`APPRam_depth*6+55)],data_in[`VWidth*(`APPRam_depth*5+56)-1:`VWidth*(`APPRam_depth*5+55)],data_in[`VWidth*(`APPRam_depth*4+56)-1:`VWidth*(`APPRam_depth*4+55)],data_in[`VWidth*(`APPRam_depth*3+56)-1:`VWidth*(`APPRam_depth*3+55)],data_in[`VWidth*(`APPRam_depth*2+56)-1:`VWidth*(`APPRam_depth*2+55)],data_in[`VWidth*(`APPRam_depth*1+56)-1:`VWidth*(`APPRam_depth*1+55)],data_in[`VWidth*(`APPRam_depth*0+56)-1:`VWidth*(`APPRam_depth*0+55)]};
			end
			56:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+57)-1:`VWidth*(`APPRam_depth*31+56)],data_in[`VWidth*(`APPRam_depth*30+57)-1:`VWidth*(`APPRam_depth*30+56)],data_in[`VWidth*(`APPRam_depth*29+57)-1:`VWidth*(`APPRam_depth*29+56)],data_in[`VWidth*(`APPRam_depth*28+57)-1:`VWidth*(`APPRam_depth*28+56)],data_in[`VWidth*(`APPRam_depth*27+57)-1:`VWidth*(`APPRam_depth*27+56)],data_in[`VWidth*(`APPRam_depth*26+57)-1:`VWidth*(`APPRam_depth*26+56)],data_in[`VWidth*(`APPRam_depth*25+57)-1:`VWidth*(`APPRam_depth*25+56)],data_in[`VWidth*(`APPRam_depth*24+57)-1:`VWidth*(`APPRam_depth*24+56)],data_in[`VWidth*(`APPRam_depth*23+57)-1:`VWidth*(`APPRam_depth*23+56)],data_in[`VWidth*(`APPRam_depth*22+57)-1:`VWidth*(`APPRam_depth*22+56)],data_in[`VWidth*(`APPRam_depth*21+57)-1:`VWidth*(`APPRam_depth*21+56)],data_in[`VWidth*(`APPRam_depth*20+57)-1:`VWidth*(`APPRam_depth*20+56)],data_in[`VWidth*(`APPRam_depth*19+57)-1:`VWidth*(`APPRam_depth*19+56)],data_in[`VWidth*(`APPRam_depth*18+57)-1:`VWidth*(`APPRam_depth*18+56)],data_in[`VWidth*(`APPRam_depth*17+57)-1:`VWidth*(`APPRam_depth*17+56)],data_in[`VWidth*(`APPRam_depth*16+57)-1:`VWidth*(`APPRam_depth*16+56)],data_in[`VWidth*(`APPRam_depth*15+57)-1:`VWidth*(`APPRam_depth*15+56)],data_in[`VWidth*(`APPRam_depth*14+57)-1:`VWidth*(`APPRam_depth*14+56)],data_in[`VWidth*(`APPRam_depth*13+57)-1:`VWidth*(`APPRam_depth*13+56)],data_in[`VWidth*(`APPRam_depth*12+57)-1:`VWidth*(`APPRam_depth*12+56)],data_in[`VWidth*(`APPRam_depth*11+57)-1:`VWidth*(`APPRam_depth*11+56)],data_in[`VWidth*(`APPRam_depth*10+57)-1:`VWidth*(`APPRam_depth*10+56)],data_in[`VWidth*(`APPRam_depth*9+57)-1:`VWidth*(`APPRam_depth*9+56)],data_in[`VWidth*(`APPRam_depth*8+57)-1:`VWidth*(`APPRam_depth*8+56)],data_in[`VWidth*(`APPRam_depth*7+57)-1:`VWidth*(`APPRam_depth*7+56)],data_in[`VWidth*(`APPRam_depth*6+57)-1:`VWidth*(`APPRam_depth*6+56)],data_in[`VWidth*(`APPRam_depth*5+57)-1:`VWidth*(`APPRam_depth*5+56)],data_in[`VWidth*(`APPRam_depth*4+57)-1:`VWidth*(`APPRam_depth*4+56)],data_in[`VWidth*(`APPRam_depth*3+57)-1:`VWidth*(`APPRam_depth*3+56)],data_in[`VWidth*(`APPRam_depth*2+57)-1:`VWidth*(`APPRam_depth*2+56)],data_in[`VWidth*(`APPRam_depth*1+57)-1:`VWidth*(`APPRam_depth*1+56)],data_in[`VWidth*(`APPRam_depth*0+57)-1:`VWidth*(`APPRam_depth*0+56)]};
			end
			57:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+58)-1:`VWidth*(`APPRam_depth*31+57)],data_in[`VWidth*(`APPRam_depth*30+58)-1:`VWidth*(`APPRam_depth*30+57)],data_in[`VWidth*(`APPRam_depth*29+58)-1:`VWidth*(`APPRam_depth*29+57)],data_in[`VWidth*(`APPRam_depth*28+58)-1:`VWidth*(`APPRam_depth*28+57)],data_in[`VWidth*(`APPRam_depth*27+58)-1:`VWidth*(`APPRam_depth*27+57)],data_in[`VWidth*(`APPRam_depth*26+58)-1:`VWidth*(`APPRam_depth*26+57)],data_in[`VWidth*(`APPRam_depth*25+58)-1:`VWidth*(`APPRam_depth*25+57)],data_in[`VWidth*(`APPRam_depth*24+58)-1:`VWidth*(`APPRam_depth*24+57)],data_in[`VWidth*(`APPRam_depth*23+58)-1:`VWidth*(`APPRam_depth*23+57)],data_in[`VWidth*(`APPRam_depth*22+58)-1:`VWidth*(`APPRam_depth*22+57)],data_in[`VWidth*(`APPRam_depth*21+58)-1:`VWidth*(`APPRam_depth*21+57)],data_in[`VWidth*(`APPRam_depth*20+58)-1:`VWidth*(`APPRam_depth*20+57)],data_in[`VWidth*(`APPRam_depth*19+58)-1:`VWidth*(`APPRam_depth*19+57)],data_in[`VWidth*(`APPRam_depth*18+58)-1:`VWidth*(`APPRam_depth*18+57)],data_in[`VWidth*(`APPRam_depth*17+58)-1:`VWidth*(`APPRam_depth*17+57)],data_in[`VWidth*(`APPRam_depth*16+58)-1:`VWidth*(`APPRam_depth*16+57)],data_in[`VWidth*(`APPRam_depth*15+58)-1:`VWidth*(`APPRam_depth*15+57)],data_in[`VWidth*(`APPRam_depth*14+58)-1:`VWidth*(`APPRam_depth*14+57)],data_in[`VWidth*(`APPRam_depth*13+58)-1:`VWidth*(`APPRam_depth*13+57)],data_in[`VWidth*(`APPRam_depth*12+58)-1:`VWidth*(`APPRam_depth*12+57)],data_in[`VWidth*(`APPRam_depth*11+58)-1:`VWidth*(`APPRam_depth*11+57)],data_in[`VWidth*(`APPRam_depth*10+58)-1:`VWidth*(`APPRam_depth*10+57)],data_in[`VWidth*(`APPRam_depth*9+58)-1:`VWidth*(`APPRam_depth*9+57)],data_in[`VWidth*(`APPRam_depth*8+58)-1:`VWidth*(`APPRam_depth*8+57)],data_in[`VWidth*(`APPRam_depth*7+58)-1:`VWidth*(`APPRam_depth*7+57)],data_in[`VWidth*(`APPRam_depth*6+58)-1:`VWidth*(`APPRam_depth*6+57)],data_in[`VWidth*(`APPRam_depth*5+58)-1:`VWidth*(`APPRam_depth*5+57)],data_in[`VWidth*(`APPRam_depth*4+58)-1:`VWidth*(`APPRam_depth*4+57)],data_in[`VWidth*(`APPRam_depth*3+58)-1:`VWidth*(`APPRam_depth*3+57)],data_in[`VWidth*(`APPRam_depth*2+58)-1:`VWidth*(`APPRam_depth*2+57)],data_in[`VWidth*(`APPRam_depth*1+58)-1:`VWidth*(`APPRam_depth*1+57)],data_in[`VWidth*(`APPRam_depth*0+58)-1:`VWidth*(`APPRam_depth*0+57)]};
			end
			58:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+59)-1:`VWidth*(`APPRam_depth*31+58)],data_in[`VWidth*(`APPRam_depth*30+59)-1:`VWidth*(`APPRam_depth*30+58)],data_in[`VWidth*(`APPRam_depth*29+59)-1:`VWidth*(`APPRam_depth*29+58)],data_in[`VWidth*(`APPRam_depth*28+59)-1:`VWidth*(`APPRam_depth*28+58)],data_in[`VWidth*(`APPRam_depth*27+59)-1:`VWidth*(`APPRam_depth*27+58)],data_in[`VWidth*(`APPRam_depth*26+59)-1:`VWidth*(`APPRam_depth*26+58)],data_in[`VWidth*(`APPRam_depth*25+59)-1:`VWidth*(`APPRam_depth*25+58)],data_in[`VWidth*(`APPRam_depth*24+59)-1:`VWidth*(`APPRam_depth*24+58)],data_in[`VWidth*(`APPRam_depth*23+59)-1:`VWidth*(`APPRam_depth*23+58)],data_in[`VWidth*(`APPRam_depth*22+59)-1:`VWidth*(`APPRam_depth*22+58)],data_in[`VWidth*(`APPRam_depth*21+59)-1:`VWidth*(`APPRam_depth*21+58)],data_in[`VWidth*(`APPRam_depth*20+59)-1:`VWidth*(`APPRam_depth*20+58)],data_in[`VWidth*(`APPRam_depth*19+59)-1:`VWidth*(`APPRam_depth*19+58)],data_in[`VWidth*(`APPRam_depth*18+59)-1:`VWidth*(`APPRam_depth*18+58)],data_in[`VWidth*(`APPRam_depth*17+59)-1:`VWidth*(`APPRam_depth*17+58)],data_in[`VWidth*(`APPRam_depth*16+59)-1:`VWidth*(`APPRam_depth*16+58)],data_in[`VWidth*(`APPRam_depth*15+59)-1:`VWidth*(`APPRam_depth*15+58)],data_in[`VWidth*(`APPRam_depth*14+59)-1:`VWidth*(`APPRam_depth*14+58)],data_in[`VWidth*(`APPRam_depth*13+59)-1:`VWidth*(`APPRam_depth*13+58)],data_in[`VWidth*(`APPRam_depth*12+59)-1:`VWidth*(`APPRam_depth*12+58)],data_in[`VWidth*(`APPRam_depth*11+59)-1:`VWidth*(`APPRam_depth*11+58)],data_in[`VWidth*(`APPRam_depth*10+59)-1:`VWidth*(`APPRam_depth*10+58)],data_in[`VWidth*(`APPRam_depth*9+59)-1:`VWidth*(`APPRam_depth*9+58)],data_in[`VWidth*(`APPRam_depth*8+59)-1:`VWidth*(`APPRam_depth*8+58)],data_in[`VWidth*(`APPRam_depth*7+59)-1:`VWidth*(`APPRam_depth*7+58)],data_in[`VWidth*(`APPRam_depth*6+59)-1:`VWidth*(`APPRam_depth*6+58)],data_in[`VWidth*(`APPRam_depth*5+59)-1:`VWidth*(`APPRam_depth*5+58)],data_in[`VWidth*(`APPRam_depth*4+59)-1:`VWidth*(`APPRam_depth*4+58)],data_in[`VWidth*(`APPRam_depth*3+59)-1:`VWidth*(`APPRam_depth*3+58)],data_in[`VWidth*(`APPRam_depth*2+59)-1:`VWidth*(`APPRam_depth*2+58)],data_in[`VWidth*(`APPRam_depth*1+59)-1:`VWidth*(`APPRam_depth*1+58)],data_in[`VWidth*(`APPRam_depth*0+59)-1:`VWidth*(`APPRam_depth*0+58)]};
			end
			59:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+60)-1:`VWidth*(`APPRam_depth*31+59)],data_in[`VWidth*(`APPRam_depth*30+60)-1:`VWidth*(`APPRam_depth*30+59)],data_in[`VWidth*(`APPRam_depth*29+60)-1:`VWidth*(`APPRam_depth*29+59)],data_in[`VWidth*(`APPRam_depth*28+60)-1:`VWidth*(`APPRam_depth*28+59)],data_in[`VWidth*(`APPRam_depth*27+60)-1:`VWidth*(`APPRam_depth*27+59)],data_in[`VWidth*(`APPRam_depth*26+60)-1:`VWidth*(`APPRam_depth*26+59)],data_in[`VWidth*(`APPRam_depth*25+60)-1:`VWidth*(`APPRam_depth*25+59)],data_in[`VWidth*(`APPRam_depth*24+60)-1:`VWidth*(`APPRam_depth*24+59)],data_in[`VWidth*(`APPRam_depth*23+60)-1:`VWidth*(`APPRam_depth*23+59)],data_in[`VWidth*(`APPRam_depth*22+60)-1:`VWidth*(`APPRam_depth*22+59)],data_in[`VWidth*(`APPRam_depth*21+60)-1:`VWidth*(`APPRam_depth*21+59)],data_in[`VWidth*(`APPRam_depth*20+60)-1:`VWidth*(`APPRam_depth*20+59)],data_in[`VWidth*(`APPRam_depth*19+60)-1:`VWidth*(`APPRam_depth*19+59)],data_in[`VWidth*(`APPRam_depth*18+60)-1:`VWidth*(`APPRam_depth*18+59)],data_in[`VWidth*(`APPRam_depth*17+60)-1:`VWidth*(`APPRam_depth*17+59)],data_in[`VWidth*(`APPRam_depth*16+60)-1:`VWidth*(`APPRam_depth*16+59)],data_in[`VWidth*(`APPRam_depth*15+60)-1:`VWidth*(`APPRam_depth*15+59)],data_in[`VWidth*(`APPRam_depth*14+60)-1:`VWidth*(`APPRam_depth*14+59)],data_in[`VWidth*(`APPRam_depth*13+60)-1:`VWidth*(`APPRam_depth*13+59)],data_in[`VWidth*(`APPRam_depth*12+60)-1:`VWidth*(`APPRam_depth*12+59)],data_in[`VWidth*(`APPRam_depth*11+60)-1:`VWidth*(`APPRam_depth*11+59)],data_in[`VWidth*(`APPRam_depth*10+60)-1:`VWidth*(`APPRam_depth*10+59)],data_in[`VWidth*(`APPRam_depth*9+60)-1:`VWidth*(`APPRam_depth*9+59)],data_in[`VWidth*(`APPRam_depth*8+60)-1:`VWidth*(`APPRam_depth*8+59)],data_in[`VWidth*(`APPRam_depth*7+60)-1:`VWidth*(`APPRam_depth*7+59)],data_in[`VWidth*(`APPRam_depth*6+60)-1:`VWidth*(`APPRam_depth*6+59)],data_in[`VWidth*(`APPRam_depth*5+60)-1:`VWidth*(`APPRam_depth*5+59)],data_in[`VWidth*(`APPRam_depth*4+60)-1:`VWidth*(`APPRam_depth*4+59)],data_in[`VWidth*(`APPRam_depth*3+60)-1:`VWidth*(`APPRam_depth*3+59)],data_in[`VWidth*(`APPRam_depth*2+60)-1:`VWidth*(`APPRam_depth*2+59)],data_in[`VWidth*(`APPRam_depth*1+60)-1:`VWidth*(`APPRam_depth*1+59)],data_in[`VWidth*(`APPRam_depth*0+60)-1:`VWidth*(`APPRam_depth*0+59)]};
			end
			60:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+61)-1:`VWidth*(`APPRam_depth*31+60)],data_in[`VWidth*(`APPRam_depth*30+61)-1:`VWidth*(`APPRam_depth*30+60)],data_in[`VWidth*(`APPRam_depth*29+61)-1:`VWidth*(`APPRam_depth*29+60)],data_in[`VWidth*(`APPRam_depth*28+61)-1:`VWidth*(`APPRam_depth*28+60)],data_in[`VWidth*(`APPRam_depth*27+61)-1:`VWidth*(`APPRam_depth*27+60)],data_in[`VWidth*(`APPRam_depth*26+61)-1:`VWidth*(`APPRam_depth*26+60)],data_in[`VWidth*(`APPRam_depth*25+61)-1:`VWidth*(`APPRam_depth*25+60)],data_in[`VWidth*(`APPRam_depth*24+61)-1:`VWidth*(`APPRam_depth*24+60)],data_in[`VWidth*(`APPRam_depth*23+61)-1:`VWidth*(`APPRam_depth*23+60)],data_in[`VWidth*(`APPRam_depth*22+61)-1:`VWidth*(`APPRam_depth*22+60)],data_in[`VWidth*(`APPRam_depth*21+61)-1:`VWidth*(`APPRam_depth*21+60)],data_in[`VWidth*(`APPRam_depth*20+61)-1:`VWidth*(`APPRam_depth*20+60)],data_in[`VWidth*(`APPRam_depth*19+61)-1:`VWidth*(`APPRam_depth*19+60)],data_in[`VWidth*(`APPRam_depth*18+61)-1:`VWidth*(`APPRam_depth*18+60)],data_in[`VWidth*(`APPRam_depth*17+61)-1:`VWidth*(`APPRam_depth*17+60)],data_in[`VWidth*(`APPRam_depth*16+61)-1:`VWidth*(`APPRam_depth*16+60)],data_in[`VWidth*(`APPRam_depth*15+61)-1:`VWidth*(`APPRam_depth*15+60)],data_in[`VWidth*(`APPRam_depth*14+61)-1:`VWidth*(`APPRam_depth*14+60)],data_in[`VWidth*(`APPRam_depth*13+61)-1:`VWidth*(`APPRam_depth*13+60)],data_in[`VWidth*(`APPRam_depth*12+61)-1:`VWidth*(`APPRam_depth*12+60)],data_in[`VWidth*(`APPRam_depth*11+61)-1:`VWidth*(`APPRam_depth*11+60)],data_in[`VWidth*(`APPRam_depth*10+61)-1:`VWidth*(`APPRam_depth*10+60)],data_in[`VWidth*(`APPRam_depth*9+61)-1:`VWidth*(`APPRam_depth*9+60)],data_in[`VWidth*(`APPRam_depth*8+61)-1:`VWidth*(`APPRam_depth*8+60)],data_in[`VWidth*(`APPRam_depth*7+61)-1:`VWidth*(`APPRam_depth*7+60)],data_in[`VWidth*(`APPRam_depth*6+61)-1:`VWidth*(`APPRam_depth*6+60)],data_in[`VWidth*(`APPRam_depth*5+61)-1:`VWidth*(`APPRam_depth*5+60)],data_in[`VWidth*(`APPRam_depth*4+61)-1:`VWidth*(`APPRam_depth*4+60)],data_in[`VWidth*(`APPRam_depth*3+61)-1:`VWidth*(`APPRam_depth*3+60)],data_in[`VWidth*(`APPRam_depth*2+61)-1:`VWidth*(`APPRam_depth*2+60)],data_in[`VWidth*(`APPRam_depth*1+61)-1:`VWidth*(`APPRam_depth*1+60)],data_in[`VWidth*(`APPRam_depth*0+61)-1:`VWidth*(`APPRam_depth*0+60)]};
			end
			61:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+62)-1:`VWidth*(`APPRam_depth*31+61)],data_in[`VWidth*(`APPRam_depth*30+62)-1:`VWidth*(`APPRam_depth*30+61)],data_in[`VWidth*(`APPRam_depth*29+62)-1:`VWidth*(`APPRam_depth*29+61)],data_in[`VWidth*(`APPRam_depth*28+62)-1:`VWidth*(`APPRam_depth*28+61)],data_in[`VWidth*(`APPRam_depth*27+62)-1:`VWidth*(`APPRam_depth*27+61)],data_in[`VWidth*(`APPRam_depth*26+62)-1:`VWidth*(`APPRam_depth*26+61)],data_in[`VWidth*(`APPRam_depth*25+62)-1:`VWidth*(`APPRam_depth*25+61)],data_in[`VWidth*(`APPRam_depth*24+62)-1:`VWidth*(`APPRam_depth*24+61)],data_in[`VWidth*(`APPRam_depth*23+62)-1:`VWidth*(`APPRam_depth*23+61)],data_in[`VWidth*(`APPRam_depth*22+62)-1:`VWidth*(`APPRam_depth*22+61)],data_in[`VWidth*(`APPRam_depth*21+62)-1:`VWidth*(`APPRam_depth*21+61)],data_in[`VWidth*(`APPRam_depth*20+62)-1:`VWidth*(`APPRam_depth*20+61)],data_in[`VWidth*(`APPRam_depth*19+62)-1:`VWidth*(`APPRam_depth*19+61)],data_in[`VWidth*(`APPRam_depth*18+62)-1:`VWidth*(`APPRam_depth*18+61)],data_in[`VWidth*(`APPRam_depth*17+62)-1:`VWidth*(`APPRam_depth*17+61)],data_in[`VWidth*(`APPRam_depth*16+62)-1:`VWidth*(`APPRam_depth*16+61)],data_in[`VWidth*(`APPRam_depth*15+62)-1:`VWidth*(`APPRam_depth*15+61)],data_in[`VWidth*(`APPRam_depth*14+62)-1:`VWidth*(`APPRam_depth*14+61)],data_in[`VWidth*(`APPRam_depth*13+62)-1:`VWidth*(`APPRam_depth*13+61)],data_in[`VWidth*(`APPRam_depth*12+62)-1:`VWidth*(`APPRam_depth*12+61)],data_in[`VWidth*(`APPRam_depth*11+62)-1:`VWidth*(`APPRam_depth*11+61)],data_in[`VWidth*(`APPRam_depth*10+62)-1:`VWidth*(`APPRam_depth*10+61)],data_in[`VWidth*(`APPRam_depth*9+62)-1:`VWidth*(`APPRam_depth*9+61)],data_in[`VWidth*(`APPRam_depth*8+62)-1:`VWidth*(`APPRam_depth*8+61)],data_in[`VWidth*(`APPRam_depth*7+62)-1:`VWidth*(`APPRam_depth*7+61)],data_in[`VWidth*(`APPRam_depth*6+62)-1:`VWidth*(`APPRam_depth*6+61)],data_in[`VWidth*(`APPRam_depth*5+62)-1:`VWidth*(`APPRam_depth*5+61)],data_in[`VWidth*(`APPRam_depth*4+62)-1:`VWidth*(`APPRam_depth*4+61)],data_in[`VWidth*(`APPRam_depth*3+62)-1:`VWidth*(`APPRam_depth*3+61)],data_in[`VWidth*(`APPRam_depth*2+62)-1:`VWidth*(`APPRam_depth*2+61)],data_in[`VWidth*(`APPRam_depth*1+62)-1:`VWidth*(`APPRam_depth*1+61)],data_in[`VWidth*(`APPRam_depth*0+62)-1:`VWidth*(`APPRam_depth*0+61)]};
			end
			62:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+63)-1:`VWidth*(`APPRam_depth*31+62)],data_in[`VWidth*(`APPRam_depth*30+63)-1:`VWidth*(`APPRam_depth*30+62)],data_in[`VWidth*(`APPRam_depth*29+63)-1:`VWidth*(`APPRam_depth*29+62)],data_in[`VWidth*(`APPRam_depth*28+63)-1:`VWidth*(`APPRam_depth*28+62)],data_in[`VWidth*(`APPRam_depth*27+63)-1:`VWidth*(`APPRam_depth*27+62)],data_in[`VWidth*(`APPRam_depth*26+63)-1:`VWidth*(`APPRam_depth*26+62)],data_in[`VWidth*(`APPRam_depth*25+63)-1:`VWidth*(`APPRam_depth*25+62)],data_in[`VWidth*(`APPRam_depth*24+63)-1:`VWidth*(`APPRam_depth*24+62)],data_in[`VWidth*(`APPRam_depth*23+63)-1:`VWidth*(`APPRam_depth*23+62)],data_in[`VWidth*(`APPRam_depth*22+63)-1:`VWidth*(`APPRam_depth*22+62)],data_in[`VWidth*(`APPRam_depth*21+63)-1:`VWidth*(`APPRam_depth*21+62)],data_in[`VWidth*(`APPRam_depth*20+63)-1:`VWidth*(`APPRam_depth*20+62)],data_in[`VWidth*(`APPRam_depth*19+63)-1:`VWidth*(`APPRam_depth*19+62)],data_in[`VWidth*(`APPRam_depth*18+63)-1:`VWidth*(`APPRam_depth*18+62)],data_in[`VWidth*(`APPRam_depth*17+63)-1:`VWidth*(`APPRam_depth*17+62)],data_in[`VWidth*(`APPRam_depth*16+63)-1:`VWidth*(`APPRam_depth*16+62)],data_in[`VWidth*(`APPRam_depth*15+63)-1:`VWidth*(`APPRam_depth*15+62)],data_in[`VWidth*(`APPRam_depth*14+63)-1:`VWidth*(`APPRam_depth*14+62)],data_in[`VWidth*(`APPRam_depth*13+63)-1:`VWidth*(`APPRam_depth*13+62)],data_in[`VWidth*(`APPRam_depth*12+63)-1:`VWidth*(`APPRam_depth*12+62)],data_in[`VWidth*(`APPRam_depth*11+63)-1:`VWidth*(`APPRam_depth*11+62)],data_in[`VWidth*(`APPRam_depth*10+63)-1:`VWidth*(`APPRam_depth*10+62)],data_in[`VWidth*(`APPRam_depth*9+63)-1:`VWidth*(`APPRam_depth*9+62)],data_in[`VWidth*(`APPRam_depth*8+63)-1:`VWidth*(`APPRam_depth*8+62)],data_in[`VWidth*(`APPRam_depth*7+63)-1:`VWidth*(`APPRam_depth*7+62)],data_in[`VWidth*(`APPRam_depth*6+63)-1:`VWidth*(`APPRam_depth*6+62)],data_in[`VWidth*(`APPRam_depth*5+63)-1:`VWidth*(`APPRam_depth*5+62)],data_in[`VWidth*(`APPRam_depth*4+63)-1:`VWidth*(`APPRam_depth*4+62)],data_in[`VWidth*(`APPRam_depth*3+63)-1:`VWidth*(`APPRam_depth*3+62)],data_in[`VWidth*(`APPRam_depth*2+63)-1:`VWidth*(`APPRam_depth*2+62)],data_in[`VWidth*(`APPRam_depth*1+63)-1:`VWidth*(`APPRam_depth*1+62)],data_in[`VWidth*(`APPRam_depth*0+63)-1:`VWidth*(`APPRam_depth*0+62)]};
			end
			63:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+64)-1:`VWidth*(`APPRam_depth*31+63)],data_in[`VWidth*(`APPRam_depth*30+64)-1:`VWidth*(`APPRam_depth*30+63)],data_in[`VWidth*(`APPRam_depth*29+64)-1:`VWidth*(`APPRam_depth*29+63)],data_in[`VWidth*(`APPRam_depth*28+64)-1:`VWidth*(`APPRam_depth*28+63)],data_in[`VWidth*(`APPRam_depth*27+64)-1:`VWidth*(`APPRam_depth*27+63)],data_in[`VWidth*(`APPRam_depth*26+64)-1:`VWidth*(`APPRam_depth*26+63)],data_in[`VWidth*(`APPRam_depth*25+64)-1:`VWidth*(`APPRam_depth*25+63)],data_in[`VWidth*(`APPRam_depth*24+64)-1:`VWidth*(`APPRam_depth*24+63)],data_in[`VWidth*(`APPRam_depth*23+64)-1:`VWidth*(`APPRam_depth*23+63)],data_in[`VWidth*(`APPRam_depth*22+64)-1:`VWidth*(`APPRam_depth*22+63)],data_in[`VWidth*(`APPRam_depth*21+64)-1:`VWidth*(`APPRam_depth*21+63)],data_in[`VWidth*(`APPRam_depth*20+64)-1:`VWidth*(`APPRam_depth*20+63)],data_in[`VWidth*(`APPRam_depth*19+64)-1:`VWidth*(`APPRam_depth*19+63)],data_in[`VWidth*(`APPRam_depth*18+64)-1:`VWidth*(`APPRam_depth*18+63)],data_in[`VWidth*(`APPRam_depth*17+64)-1:`VWidth*(`APPRam_depth*17+63)],data_in[`VWidth*(`APPRam_depth*16+64)-1:`VWidth*(`APPRam_depth*16+63)],data_in[`VWidth*(`APPRam_depth*15+64)-1:`VWidth*(`APPRam_depth*15+63)],data_in[`VWidth*(`APPRam_depth*14+64)-1:`VWidth*(`APPRam_depth*14+63)],data_in[`VWidth*(`APPRam_depth*13+64)-1:`VWidth*(`APPRam_depth*13+63)],data_in[`VWidth*(`APPRam_depth*12+64)-1:`VWidth*(`APPRam_depth*12+63)],data_in[`VWidth*(`APPRam_depth*11+64)-1:`VWidth*(`APPRam_depth*11+63)],data_in[`VWidth*(`APPRam_depth*10+64)-1:`VWidth*(`APPRam_depth*10+63)],data_in[`VWidth*(`APPRam_depth*9+64)-1:`VWidth*(`APPRam_depth*9+63)],data_in[`VWidth*(`APPRam_depth*8+64)-1:`VWidth*(`APPRam_depth*8+63)],data_in[`VWidth*(`APPRam_depth*7+64)-1:`VWidth*(`APPRam_depth*7+63)],data_in[`VWidth*(`APPRam_depth*6+64)-1:`VWidth*(`APPRam_depth*6+63)],data_in[`VWidth*(`APPRam_depth*5+64)-1:`VWidth*(`APPRam_depth*5+63)],data_in[`VWidth*(`APPRam_depth*4+64)-1:`VWidth*(`APPRam_depth*4+63)],data_in[`VWidth*(`APPRam_depth*3+64)-1:`VWidth*(`APPRam_depth*3+63)],data_in[`VWidth*(`APPRam_depth*2+64)-1:`VWidth*(`APPRam_depth*2+63)],data_in[`VWidth*(`APPRam_depth*1+64)-1:`VWidth*(`APPRam_depth*1+63)],data_in[`VWidth*(`APPRam_depth*0+64)-1:`VWidth*(`APPRam_depth*0+63)]};
			end
			64:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+65)-1:`VWidth*(`APPRam_depth*31+64)],data_in[`VWidth*(`APPRam_depth*30+65)-1:`VWidth*(`APPRam_depth*30+64)],data_in[`VWidth*(`APPRam_depth*29+65)-1:`VWidth*(`APPRam_depth*29+64)],data_in[`VWidth*(`APPRam_depth*28+65)-1:`VWidth*(`APPRam_depth*28+64)],data_in[`VWidth*(`APPRam_depth*27+65)-1:`VWidth*(`APPRam_depth*27+64)],data_in[`VWidth*(`APPRam_depth*26+65)-1:`VWidth*(`APPRam_depth*26+64)],data_in[`VWidth*(`APPRam_depth*25+65)-1:`VWidth*(`APPRam_depth*25+64)],data_in[`VWidth*(`APPRam_depth*24+65)-1:`VWidth*(`APPRam_depth*24+64)],data_in[`VWidth*(`APPRam_depth*23+65)-1:`VWidth*(`APPRam_depth*23+64)],data_in[`VWidth*(`APPRam_depth*22+65)-1:`VWidth*(`APPRam_depth*22+64)],data_in[`VWidth*(`APPRam_depth*21+65)-1:`VWidth*(`APPRam_depth*21+64)],data_in[`VWidth*(`APPRam_depth*20+65)-1:`VWidth*(`APPRam_depth*20+64)],data_in[`VWidth*(`APPRam_depth*19+65)-1:`VWidth*(`APPRam_depth*19+64)],data_in[`VWidth*(`APPRam_depth*18+65)-1:`VWidth*(`APPRam_depth*18+64)],data_in[`VWidth*(`APPRam_depth*17+65)-1:`VWidth*(`APPRam_depth*17+64)],data_in[`VWidth*(`APPRam_depth*16+65)-1:`VWidth*(`APPRam_depth*16+64)],data_in[`VWidth*(`APPRam_depth*15+65)-1:`VWidth*(`APPRam_depth*15+64)],data_in[`VWidth*(`APPRam_depth*14+65)-1:`VWidth*(`APPRam_depth*14+64)],data_in[`VWidth*(`APPRam_depth*13+65)-1:`VWidth*(`APPRam_depth*13+64)],data_in[`VWidth*(`APPRam_depth*12+65)-1:`VWidth*(`APPRam_depth*12+64)],data_in[`VWidth*(`APPRam_depth*11+65)-1:`VWidth*(`APPRam_depth*11+64)],data_in[`VWidth*(`APPRam_depth*10+65)-1:`VWidth*(`APPRam_depth*10+64)],data_in[`VWidth*(`APPRam_depth*9+65)-1:`VWidth*(`APPRam_depth*9+64)],data_in[`VWidth*(`APPRam_depth*8+65)-1:`VWidth*(`APPRam_depth*8+64)],data_in[`VWidth*(`APPRam_depth*7+65)-1:`VWidth*(`APPRam_depth*7+64)],data_in[`VWidth*(`APPRam_depth*6+65)-1:`VWidth*(`APPRam_depth*6+64)],data_in[`VWidth*(`APPRam_depth*5+65)-1:`VWidth*(`APPRam_depth*5+64)],data_in[`VWidth*(`APPRam_depth*4+65)-1:`VWidth*(`APPRam_depth*4+64)],data_in[`VWidth*(`APPRam_depth*3+65)-1:`VWidth*(`APPRam_depth*3+64)],data_in[`VWidth*(`APPRam_depth*2+65)-1:`VWidth*(`APPRam_depth*2+64)],data_in[`VWidth*(`APPRam_depth*1+65)-1:`VWidth*(`APPRam_depth*1+64)],data_in[`VWidth*(`APPRam_depth*0+65)-1:`VWidth*(`APPRam_depth*0+64)]};
			end
			65:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+66)-1:`VWidth*(`APPRam_depth*31+65)],data_in[`VWidth*(`APPRam_depth*30+66)-1:`VWidth*(`APPRam_depth*30+65)],data_in[`VWidth*(`APPRam_depth*29+66)-1:`VWidth*(`APPRam_depth*29+65)],data_in[`VWidth*(`APPRam_depth*28+66)-1:`VWidth*(`APPRam_depth*28+65)],data_in[`VWidth*(`APPRam_depth*27+66)-1:`VWidth*(`APPRam_depth*27+65)],data_in[`VWidth*(`APPRam_depth*26+66)-1:`VWidth*(`APPRam_depth*26+65)],data_in[`VWidth*(`APPRam_depth*25+66)-1:`VWidth*(`APPRam_depth*25+65)],data_in[`VWidth*(`APPRam_depth*24+66)-1:`VWidth*(`APPRam_depth*24+65)],data_in[`VWidth*(`APPRam_depth*23+66)-1:`VWidth*(`APPRam_depth*23+65)],data_in[`VWidth*(`APPRam_depth*22+66)-1:`VWidth*(`APPRam_depth*22+65)],data_in[`VWidth*(`APPRam_depth*21+66)-1:`VWidth*(`APPRam_depth*21+65)],data_in[`VWidth*(`APPRam_depth*20+66)-1:`VWidth*(`APPRam_depth*20+65)],data_in[`VWidth*(`APPRam_depth*19+66)-1:`VWidth*(`APPRam_depth*19+65)],data_in[`VWidth*(`APPRam_depth*18+66)-1:`VWidth*(`APPRam_depth*18+65)],data_in[`VWidth*(`APPRam_depth*17+66)-1:`VWidth*(`APPRam_depth*17+65)],data_in[`VWidth*(`APPRam_depth*16+66)-1:`VWidth*(`APPRam_depth*16+65)],data_in[`VWidth*(`APPRam_depth*15+66)-1:`VWidth*(`APPRam_depth*15+65)],data_in[`VWidth*(`APPRam_depth*14+66)-1:`VWidth*(`APPRam_depth*14+65)],data_in[`VWidth*(`APPRam_depth*13+66)-1:`VWidth*(`APPRam_depth*13+65)],data_in[`VWidth*(`APPRam_depth*12+66)-1:`VWidth*(`APPRam_depth*12+65)],data_in[`VWidth*(`APPRam_depth*11+66)-1:`VWidth*(`APPRam_depth*11+65)],data_in[`VWidth*(`APPRam_depth*10+66)-1:`VWidth*(`APPRam_depth*10+65)],data_in[`VWidth*(`APPRam_depth*9+66)-1:`VWidth*(`APPRam_depth*9+65)],data_in[`VWidth*(`APPRam_depth*8+66)-1:`VWidth*(`APPRam_depth*8+65)],data_in[`VWidth*(`APPRam_depth*7+66)-1:`VWidth*(`APPRam_depth*7+65)],data_in[`VWidth*(`APPRam_depth*6+66)-1:`VWidth*(`APPRam_depth*6+65)],data_in[`VWidth*(`APPRam_depth*5+66)-1:`VWidth*(`APPRam_depth*5+65)],data_in[`VWidth*(`APPRam_depth*4+66)-1:`VWidth*(`APPRam_depth*4+65)],data_in[`VWidth*(`APPRam_depth*3+66)-1:`VWidth*(`APPRam_depth*3+65)],data_in[`VWidth*(`APPRam_depth*2+66)-1:`VWidth*(`APPRam_depth*2+65)],data_in[`VWidth*(`APPRam_depth*1+66)-1:`VWidth*(`APPRam_depth*1+65)],data_in[`VWidth*(`APPRam_depth*0+66)-1:`VWidth*(`APPRam_depth*0+65)]};
			end
			66:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+67)-1:`VWidth*(`APPRam_depth*31+66)],data_in[`VWidth*(`APPRam_depth*30+67)-1:`VWidth*(`APPRam_depth*30+66)],data_in[`VWidth*(`APPRam_depth*29+67)-1:`VWidth*(`APPRam_depth*29+66)],data_in[`VWidth*(`APPRam_depth*28+67)-1:`VWidth*(`APPRam_depth*28+66)],data_in[`VWidth*(`APPRam_depth*27+67)-1:`VWidth*(`APPRam_depth*27+66)],data_in[`VWidth*(`APPRam_depth*26+67)-1:`VWidth*(`APPRam_depth*26+66)],data_in[`VWidth*(`APPRam_depth*25+67)-1:`VWidth*(`APPRam_depth*25+66)],data_in[`VWidth*(`APPRam_depth*24+67)-1:`VWidth*(`APPRam_depth*24+66)],data_in[`VWidth*(`APPRam_depth*23+67)-1:`VWidth*(`APPRam_depth*23+66)],data_in[`VWidth*(`APPRam_depth*22+67)-1:`VWidth*(`APPRam_depth*22+66)],data_in[`VWidth*(`APPRam_depth*21+67)-1:`VWidth*(`APPRam_depth*21+66)],data_in[`VWidth*(`APPRam_depth*20+67)-1:`VWidth*(`APPRam_depth*20+66)],data_in[`VWidth*(`APPRam_depth*19+67)-1:`VWidth*(`APPRam_depth*19+66)],data_in[`VWidth*(`APPRam_depth*18+67)-1:`VWidth*(`APPRam_depth*18+66)],data_in[`VWidth*(`APPRam_depth*17+67)-1:`VWidth*(`APPRam_depth*17+66)],data_in[`VWidth*(`APPRam_depth*16+67)-1:`VWidth*(`APPRam_depth*16+66)],data_in[`VWidth*(`APPRam_depth*15+67)-1:`VWidth*(`APPRam_depth*15+66)],data_in[`VWidth*(`APPRam_depth*14+67)-1:`VWidth*(`APPRam_depth*14+66)],data_in[`VWidth*(`APPRam_depth*13+67)-1:`VWidth*(`APPRam_depth*13+66)],data_in[`VWidth*(`APPRam_depth*12+67)-1:`VWidth*(`APPRam_depth*12+66)],data_in[`VWidth*(`APPRam_depth*11+67)-1:`VWidth*(`APPRam_depth*11+66)],data_in[`VWidth*(`APPRam_depth*10+67)-1:`VWidth*(`APPRam_depth*10+66)],data_in[`VWidth*(`APPRam_depth*9+67)-1:`VWidth*(`APPRam_depth*9+66)],data_in[`VWidth*(`APPRam_depth*8+67)-1:`VWidth*(`APPRam_depth*8+66)],data_in[`VWidth*(`APPRam_depth*7+67)-1:`VWidth*(`APPRam_depth*7+66)],data_in[`VWidth*(`APPRam_depth*6+67)-1:`VWidth*(`APPRam_depth*6+66)],data_in[`VWidth*(`APPRam_depth*5+67)-1:`VWidth*(`APPRam_depth*5+66)],data_in[`VWidth*(`APPRam_depth*4+67)-1:`VWidth*(`APPRam_depth*4+66)],data_in[`VWidth*(`APPRam_depth*3+67)-1:`VWidth*(`APPRam_depth*3+66)],data_in[`VWidth*(`APPRam_depth*2+67)-1:`VWidth*(`APPRam_depth*2+66)],data_in[`VWidth*(`APPRam_depth*1+67)-1:`VWidth*(`APPRam_depth*1+66)],data_in[`VWidth*(`APPRam_depth*0+67)-1:`VWidth*(`APPRam_depth*0+66)]};
			end
			67:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+68)-1:`VWidth*(`APPRam_depth*31+67)],data_in[`VWidth*(`APPRam_depth*30+68)-1:`VWidth*(`APPRam_depth*30+67)],data_in[`VWidth*(`APPRam_depth*29+68)-1:`VWidth*(`APPRam_depth*29+67)],data_in[`VWidth*(`APPRam_depth*28+68)-1:`VWidth*(`APPRam_depth*28+67)],data_in[`VWidth*(`APPRam_depth*27+68)-1:`VWidth*(`APPRam_depth*27+67)],data_in[`VWidth*(`APPRam_depth*26+68)-1:`VWidth*(`APPRam_depth*26+67)],data_in[`VWidth*(`APPRam_depth*25+68)-1:`VWidth*(`APPRam_depth*25+67)],data_in[`VWidth*(`APPRam_depth*24+68)-1:`VWidth*(`APPRam_depth*24+67)],data_in[`VWidth*(`APPRam_depth*23+68)-1:`VWidth*(`APPRam_depth*23+67)],data_in[`VWidth*(`APPRam_depth*22+68)-1:`VWidth*(`APPRam_depth*22+67)],data_in[`VWidth*(`APPRam_depth*21+68)-1:`VWidth*(`APPRam_depth*21+67)],data_in[`VWidth*(`APPRam_depth*20+68)-1:`VWidth*(`APPRam_depth*20+67)],data_in[`VWidth*(`APPRam_depth*19+68)-1:`VWidth*(`APPRam_depth*19+67)],data_in[`VWidth*(`APPRam_depth*18+68)-1:`VWidth*(`APPRam_depth*18+67)],data_in[`VWidth*(`APPRam_depth*17+68)-1:`VWidth*(`APPRam_depth*17+67)],data_in[`VWidth*(`APPRam_depth*16+68)-1:`VWidth*(`APPRam_depth*16+67)],data_in[`VWidth*(`APPRam_depth*15+68)-1:`VWidth*(`APPRam_depth*15+67)],data_in[`VWidth*(`APPRam_depth*14+68)-1:`VWidth*(`APPRam_depth*14+67)],data_in[`VWidth*(`APPRam_depth*13+68)-1:`VWidth*(`APPRam_depth*13+67)],data_in[`VWidth*(`APPRam_depth*12+68)-1:`VWidth*(`APPRam_depth*12+67)],data_in[`VWidth*(`APPRam_depth*11+68)-1:`VWidth*(`APPRam_depth*11+67)],data_in[`VWidth*(`APPRam_depth*10+68)-1:`VWidth*(`APPRam_depth*10+67)],data_in[`VWidth*(`APPRam_depth*9+68)-1:`VWidth*(`APPRam_depth*9+67)],data_in[`VWidth*(`APPRam_depth*8+68)-1:`VWidth*(`APPRam_depth*8+67)],data_in[`VWidth*(`APPRam_depth*7+68)-1:`VWidth*(`APPRam_depth*7+67)],data_in[`VWidth*(`APPRam_depth*6+68)-1:`VWidth*(`APPRam_depth*6+67)],data_in[`VWidth*(`APPRam_depth*5+68)-1:`VWidth*(`APPRam_depth*5+67)],data_in[`VWidth*(`APPRam_depth*4+68)-1:`VWidth*(`APPRam_depth*4+67)],data_in[`VWidth*(`APPRam_depth*3+68)-1:`VWidth*(`APPRam_depth*3+67)],data_in[`VWidth*(`APPRam_depth*2+68)-1:`VWidth*(`APPRam_depth*2+67)],data_in[`VWidth*(`APPRam_depth*1+68)-1:`VWidth*(`APPRam_depth*1+67)],data_in[`VWidth*(`APPRam_depth*0+68)-1:`VWidth*(`APPRam_depth*0+67)]};
			end
			68:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+69)-1:`VWidth*(`APPRam_depth*31+68)],data_in[`VWidth*(`APPRam_depth*30+69)-1:`VWidth*(`APPRam_depth*30+68)],data_in[`VWidth*(`APPRam_depth*29+69)-1:`VWidth*(`APPRam_depth*29+68)],data_in[`VWidth*(`APPRam_depth*28+69)-1:`VWidth*(`APPRam_depth*28+68)],data_in[`VWidth*(`APPRam_depth*27+69)-1:`VWidth*(`APPRam_depth*27+68)],data_in[`VWidth*(`APPRam_depth*26+69)-1:`VWidth*(`APPRam_depth*26+68)],data_in[`VWidth*(`APPRam_depth*25+69)-1:`VWidth*(`APPRam_depth*25+68)],data_in[`VWidth*(`APPRam_depth*24+69)-1:`VWidth*(`APPRam_depth*24+68)],data_in[`VWidth*(`APPRam_depth*23+69)-1:`VWidth*(`APPRam_depth*23+68)],data_in[`VWidth*(`APPRam_depth*22+69)-1:`VWidth*(`APPRam_depth*22+68)],data_in[`VWidth*(`APPRam_depth*21+69)-1:`VWidth*(`APPRam_depth*21+68)],data_in[`VWidth*(`APPRam_depth*20+69)-1:`VWidth*(`APPRam_depth*20+68)],data_in[`VWidth*(`APPRam_depth*19+69)-1:`VWidth*(`APPRam_depth*19+68)],data_in[`VWidth*(`APPRam_depth*18+69)-1:`VWidth*(`APPRam_depth*18+68)],data_in[`VWidth*(`APPRam_depth*17+69)-1:`VWidth*(`APPRam_depth*17+68)],data_in[`VWidth*(`APPRam_depth*16+69)-1:`VWidth*(`APPRam_depth*16+68)],data_in[`VWidth*(`APPRam_depth*15+69)-1:`VWidth*(`APPRam_depth*15+68)],data_in[`VWidth*(`APPRam_depth*14+69)-1:`VWidth*(`APPRam_depth*14+68)],data_in[`VWidth*(`APPRam_depth*13+69)-1:`VWidth*(`APPRam_depth*13+68)],data_in[`VWidth*(`APPRam_depth*12+69)-1:`VWidth*(`APPRam_depth*12+68)],data_in[`VWidth*(`APPRam_depth*11+69)-1:`VWidth*(`APPRam_depth*11+68)],data_in[`VWidth*(`APPRam_depth*10+69)-1:`VWidth*(`APPRam_depth*10+68)],data_in[`VWidth*(`APPRam_depth*9+69)-1:`VWidth*(`APPRam_depth*9+68)],data_in[`VWidth*(`APPRam_depth*8+69)-1:`VWidth*(`APPRam_depth*8+68)],data_in[`VWidth*(`APPRam_depth*7+69)-1:`VWidth*(`APPRam_depth*7+68)],data_in[`VWidth*(`APPRam_depth*6+69)-1:`VWidth*(`APPRam_depth*6+68)],data_in[`VWidth*(`APPRam_depth*5+69)-1:`VWidth*(`APPRam_depth*5+68)],data_in[`VWidth*(`APPRam_depth*4+69)-1:`VWidth*(`APPRam_depth*4+68)],data_in[`VWidth*(`APPRam_depth*3+69)-1:`VWidth*(`APPRam_depth*3+68)],data_in[`VWidth*(`APPRam_depth*2+69)-1:`VWidth*(`APPRam_depth*2+68)],data_in[`VWidth*(`APPRam_depth*1+69)-1:`VWidth*(`APPRam_depth*1+68)],data_in[`VWidth*(`APPRam_depth*0+69)-1:`VWidth*(`APPRam_depth*0+68)]};
			end
			69:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+70)-1:`VWidth*(`APPRam_depth*31+69)],data_in[`VWidth*(`APPRam_depth*30+70)-1:`VWidth*(`APPRam_depth*30+69)],data_in[`VWidth*(`APPRam_depth*29+70)-1:`VWidth*(`APPRam_depth*29+69)],data_in[`VWidth*(`APPRam_depth*28+70)-1:`VWidth*(`APPRam_depth*28+69)],data_in[`VWidth*(`APPRam_depth*27+70)-1:`VWidth*(`APPRam_depth*27+69)],data_in[`VWidth*(`APPRam_depth*26+70)-1:`VWidth*(`APPRam_depth*26+69)],data_in[`VWidth*(`APPRam_depth*25+70)-1:`VWidth*(`APPRam_depth*25+69)],data_in[`VWidth*(`APPRam_depth*24+70)-1:`VWidth*(`APPRam_depth*24+69)],data_in[`VWidth*(`APPRam_depth*23+70)-1:`VWidth*(`APPRam_depth*23+69)],data_in[`VWidth*(`APPRam_depth*22+70)-1:`VWidth*(`APPRam_depth*22+69)],data_in[`VWidth*(`APPRam_depth*21+70)-1:`VWidth*(`APPRam_depth*21+69)],data_in[`VWidth*(`APPRam_depth*20+70)-1:`VWidth*(`APPRam_depth*20+69)],data_in[`VWidth*(`APPRam_depth*19+70)-1:`VWidth*(`APPRam_depth*19+69)],data_in[`VWidth*(`APPRam_depth*18+70)-1:`VWidth*(`APPRam_depth*18+69)],data_in[`VWidth*(`APPRam_depth*17+70)-1:`VWidth*(`APPRam_depth*17+69)],data_in[`VWidth*(`APPRam_depth*16+70)-1:`VWidth*(`APPRam_depth*16+69)],data_in[`VWidth*(`APPRam_depth*15+70)-1:`VWidth*(`APPRam_depth*15+69)],data_in[`VWidth*(`APPRam_depth*14+70)-1:`VWidth*(`APPRam_depth*14+69)],data_in[`VWidth*(`APPRam_depth*13+70)-1:`VWidth*(`APPRam_depth*13+69)],data_in[`VWidth*(`APPRam_depth*12+70)-1:`VWidth*(`APPRam_depth*12+69)],data_in[`VWidth*(`APPRam_depth*11+70)-1:`VWidth*(`APPRam_depth*11+69)],data_in[`VWidth*(`APPRam_depth*10+70)-1:`VWidth*(`APPRam_depth*10+69)],data_in[`VWidth*(`APPRam_depth*9+70)-1:`VWidth*(`APPRam_depth*9+69)],data_in[`VWidth*(`APPRam_depth*8+70)-1:`VWidth*(`APPRam_depth*8+69)],data_in[`VWidth*(`APPRam_depth*7+70)-1:`VWidth*(`APPRam_depth*7+69)],data_in[`VWidth*(`APPRam_depth*6+70)-1:`VWidth*(`APPRam_depth*6+69)],data_in[`VWidth*(`APPRam_depth*5+70)-1:`VWidth*(`APPRam_depth*5+69)],data_in[`VWidth*(`APPRam_depth*4+70)-1:`VWidth*(`APPRam_depth*4+69)],data_in[`VWidth*(`APPRam_depth*3+70)-1:`VWidth*(`APPRam_depth*3+69)],data_in[`VWidth*(`APPRam_depth*2+70)-1:`VWidth*(`APPRam_depth*2+69)],data_in[`VWidth*(`APPRam_depth*1+70)-1:`VWidth*(`APPRam_depth*1+69)],data_in[`VWidth*(`APPRam_depth*0+70)-1:`VWidth*(`APPRam_depth*0+69)]};
			end
			70:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+71)-1:`VWidth*(`APPRam_depth*31+70)],data_in[`VWidth*(`APPRam_depth*30+71)-1:`VWidth*(`APPRam_depth*30+70)],data_in[`VWidth*(`APPRam_depth*29+71)-1:`VWidth*(`APPRam_depth*29+70)],data_in[`VWidth*(`APPRam_depth*28+71)-1:`VWidth*(`APPRam_depth*28+70)],data_in[`VWidth*(`APPRam_depth*27+71)-1:`VWidth*(`APPRam_depth*27+70)],data_in[`VWidth*(`APPRam_depth*26+71)-1:`VWidth*(`APPRam_depth*26+70)],data_in[`VWidth*(`APPRam_depth*25+71)-1:`VWidth*(`APPRam_depth*25+70)],data_in[`VWidth*(`APPRam_depth*24+71)-1:`VWidth*(`APPRam_depth*24+70)],data_in[`VWidth*(`APPRam_depth*23+71)-1:`VWidth*(`APPRam_depth*23+70)],data_in[`VWidth*(`APPRam_depth*22+71)-1:`VWidth*(`APPRam_depth*22+70)],data_in[`VWidth*(`APPRam_depth*21+71)-1:`VWidth*(`APPRam_depth*21+70)],data_in[`VWidth*(`APPRam_depth*20+71)-1:`VWidth*(`APPRam_depth*20+70)],data_in[`VWidth*(`APPRam_depth*19+71)-1:`VWidth*(`APPRam_depth*19+70)],data_in[`VWidth*(`APPRam_depth*18+71)-1:`VWidth*(`APPRam_depth*18+70)],data_in[`VWidth*(`APPRam_depth*17+71)-1:`VWidth*(`APPRam_depth*17+70)],data_in[`VWidth*(`APPRam_depth*16+71)-1:`VWidth*(`APPRam_depth*16+70)],data_in[`VWidth*(`APPRam_depth*15+71)-1:`VWidth*(`APPRam_depth*15+70)],data_in[`VWidth*(`APPRam_depth*14+71)-1:`VWidth*(`APPRam_depth*14+70)],data_in[`VWidth*(`APPRam_depth*13+71)-1:`VWidth*(`APPRam_depth*13+70)],data_in[`VWidth*(`APPRam_depth*12+71)-1:`VWidth*(`APPRam_depth*12+70)],data_in[`VWidth*(`APPRam_depth*11+71)-1:`VWidth*(`APPRam_depth*11+70)],data_in[`VWidth*(`APPRam_depth*10+71)-1:`VWidth*(`APPRam_depth*10+70)],data_in[`VWidth*(`APPRam_depth*9+71)-1:`VWidth*(`APPRam_depth*9+70)],data_in[`VWidth*(`APPRam_depth*8+71)-1:`VWidth*(`APPRam_depth*8+70)],data_in[`VWidth*(`APPRam_depth*7+71)-1:`VWidth*(`APPRam_depth*7+70)],data_in[`VWidth*(`APPRam_depth*6+71)-1:`VWidth*(`APPRam_depth*6+70)],data_in[`VWidth*(`APPRam_depth*5+71)-1:`VWidth*(`APPRam_depth*5+70)],data_in[`VWidth*(`APPRam_depth*4+71)-1:`VWidth*(`APPRam_depth*4+70)],data_in[`VWidth*(`APPRam_depth*3+71)-1:`VWidth*(`APPRam_depth*3+70)],data_in[`VWidth*(`APPRam_depth*2+71)-1:`VWidth*(`APPRam_depth*2+70)],data_in[`VWidth*(`APPRam_depth*1+71)-1:`VWidth*(`APPRam_depth*1+70)],data_in[`VWidth*(`APPRam_depth*0+71)-1:`VWidth*(`APPRam_depth*0+70)]};
			end
			71:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+72)-1:`VWidth*(`APPRam_depth*31+71)],data_in[`VWidth*(`APPRam_depth*30+72)-1:`VWidth*(`APPRam_depth*30+71)],data_in[`VWidth*(`APPRam_depth*29+72)-1:`VWidth*(`APPRam_depth*29+71)],data_in[`VWidth*(`APPRam_depth*28+72)-1:`VWidth*(`APPRam_depth*28+71)],data_in[`VWidth*(`APPRam_depth*27+72)-1:`VWidth*(`APPRam_depth*27+71)],data_in[`VWidth*(`APPRam_depth*26+72)-1:`VWidth*(`APPRam_depth*26+71)],data_in[`VWidth*(`APPRam_depth*25+72)-1:`VWidth*(`APPRam_depth*25+71)],data_in[`VWidth*(`APPRam_depth*24+72)-1:`VWidth*(`APPRam_depth*24+71)],data_in[`VWidth*(`APPRam_depth*23+72)-1:`VWidth*(`APPRam_depth*23+71)],data_in[`VWidth*(`APPRam_depth*22+72)-1:`VWidth*(`APPRam_depth*22+71)],data_in[`VWidth*(`APPRam_depth*21+72)-1:`VWidth*(`APPRam_depth*21+71)],data_in[`VWidth*(`APPRam_depth*20+72)-1:`VWidth*(`APPRam_depth*20+71)],data_in[`VWidth*(`APPRam_depth*19+72)-1:`VWidth*(`APPRam_depth*19+71)],data_in[`VWidth*(`APPRam_depth*18+72)-1:`VWidth*(`APPRam_depth*18+71)],data_in[`VWidth*(`APPRam_depth*17+72)-1:`VWidth*(`APPRam_depth*17+71)],data_in[`VWidth*(`APPRam_depth*16+72)-1:`VWidth*(`APPRam_depth*16+71)],data_in[`VWidth*(`APPRam_depth*15+72)-1:`VWidth*(`APPRam_depth*15+71)],data_in[`VWidth*(`APPRam_depth*14+72)-1:`VWidth*(`APPRam_depth*14+71)],data_in[`VWidth*(`APPRam_depth*13+72)-1:`VWidth*(`APPRam_depth*13+71)],data_in[`VWidth*(`APPRam_depth*12+72)-1:`VWidth*(`APPRam_depth*12+71)],data_in[`VWidth*(`APPRam_depth*11+72)-1:`VWidth*(`APPRam_depth*11+71)],data_in[`VWidth*(`APPRam_depth*10+72)-1:`VWidth*(`APPRam_depth*10+71)],data_in[`VWidth*(`APPRam_depth*9+72)-1:`VWidth*(`APPRam_depth*9+71)],data_in[`VWidth*(`APPRam_depth*8+72)-1:`VWidth*(`APPRam_depth*8+71)],data_in[`VWidth*(`APPRam_depth*7+72)-1:`VWidth*(`APPRam_depth*7+71)],data_in[`VWidth*(`APPRam_depth*6+72)-1:`VWidth*(`APPRam_depth*6+71)],data_in[`VWidth*(`APPRam_depth*5+72)-1:`VWidth*(`APPRam_depth*5+71)],data_in[`VWidth*(`APPRam_depth*4+72)-1:`VWidth*(`APPRam_depth*4+71)],data_in[`VWidth*(`APPRam_depth*3+72)-1:`VWidth*(`APPRam_depth*3+71)],data_in[`VWidth*(`APPRam_depth*2+72)-1:`VWidth*(`APPRam_depth*2+71)],data_in[`VWidth*(`APPRam_depth*1+72)-1:`VWidth*(`APPRam_depth*1+71)],data_in[`VWidth*(`APPRam_depth*0+72)-1:`VWidth*(`APPRam_depth*0+71)]};
			end
			72:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+73)-1:`VWidth*(`APPRam_depth*31+72)],data_in[`VWidth*(`APPRam_depth*30+73)-1:`VWidth*(`APPRam_depth*30+72)],data_in[`VWidth*(`APPRam_depth*29+73)-1:`VWidth*(`APPRam_depth*29+72)],data_in[`VWidth*(`APPRam_depth*28+73)-1:`VWidth*(`APPRam_depth*28+72)],data_in[`VWidth*(`APPRam_depth*27+73)-1:`VWidth*(`APPRam_depth*27+72)],data_in[`VWidth*(`APPRam_depth*26+73)-1:`VWidth*(`APPRam_depth*26+72)],data_in[`VWidth*(`APPRam_depth*25+73)-1:`VWidth*(`APPRam_depth*25+72)],data_in[`VWidth*(`APPRam_depth*24+73)-1:`VWidth*(`APPRam_depth*24+72)],data_in[`VWidth*(`APPRam_depth*23+73)-1:`VWidth*(`APPRam_depth*23+72)],data_in[`VWidth*(`APPRam_depth*22+73)-1:`VWidth*(`APPRam_depth*22+72)],data_in[`VWidth*(`APPRam_depth*21+73)-1:`VWidth*(`APPRam_depth*21+72)],data_in[`VWidth*(`APPRam_depth*20+73)-1:`VWidth*(`APPRam_depth*20+72)],data_in[`VWidth*(`APPRam_depth*19+73)-1:`VWidth*(`APPRam_depth*19+72)],data_in[`VWidth*(`APPRam_depth*18+73)-1:`VWidth*(`APPRam_depth*18+72)],data_in[`VWidth*(`APPRam_depth*17+73)-1:`VWidth*(`APPRam_depth*17+72)],data_in[`VWidth*(`APPRam_depth*16+73)-1:`VWidth*(`APPRam_depth*16+72)],data_in[`VWidth*(`APPRam_depth*15+73)-1:`VWidth*(`APPRam_depth*15+72)],data_in[`VWidth*(`APPRam_depth*14+73)-1:`VWidth*(`APPRam_depth*14+72)],data_in[`VWidth*(`APPRam_depth*13+73)-1:`VWidth*(`APPRam_depth*13+72)],data_in[`VWidth*(`APPRam_depth*12+73)-1:`VWidth*(`APPRam_depth*12+72)],data_in[`VWidth*(`APPRam_depth*11+73)-1:`VWidth*(`APPRam_depth*11+72)],data_in[`VWidth*(`APPRam_depth*10+73)-1:`VWidth*(`APPRam_depth*10+72)],data_in[`VWidth*(`APPRam_depth*9+73)-1:`VWidth*(`APPRam_depth*9+72)],data_in[`VWidth*(`APPRam_depth*8+73)-1:`VWidth*(`APPRam_depth*8+72)],data_in[`VWidth*(`APPRam_depth*7+73)-1:`VWidth*(`APPRam_depth*7+72)],data_in[`VWidth*(`APPRam_depth*6+73)-1:`VWidth*(`APPRam_depth*6+72)],data_in[`VWidth*(`APPRam_depth*5+73)-1:`VWidth*(`APPRam_depth*5+72)],data_in[`VWidth*(`APPRam_depth*4+73)-1:`VWidth*(`APPRam_depth*4+72)],data_in[`VWidth*(`APPRam_depth*3+73)-1:`VWidth*(`APPRam_depth*3+72)],data_in[`VWidth*(`APPRam_depth*2+73)-1:`VWidth*(`APPRam_depth*2+72)],data_in[`VWidth*(`APPRam_depth*1+73)-1:`VWidth*(`APPRam_depth*1+72)],data_in[`VWidth*(`APPRam_depth*0+73)-1:`VWidth*(`APPRam_depth*0+72)]};
			end
			73:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+74)-1:`VWidth*(`APPRam_depth*31+73)],data_in[`VWidth*(`APPRam_depth*30+74)-1:`VWidth*(`APPRam_depth*30+73)],data_in[`VWidth*(`APPRam_depth*29+74)-1:`VWidth*(`APPRam_depth*29+73)],data_in[`VWidth*(`APPRam_depth*28+74)-1:`VWidth*(`APPRam_depth*28+73)],data_in[`VWidth*(`APPRam_depth*27+74)-1:`VWidth*(`APPRam_depth*27+73)],data_in[`VWidth*(`APPRam_depth*26+74)-1:`VWidth*(`APPRam_depth*26+73)],data_in[`VWidth*(`APPRam_depth*25+74)-1:`VWidth*(`APPRam_depth*25+73)],data_in[`VWidth*(`APPRam_depth*24+74)-1:`VWidth*(`APPRam_depth*24+73)],data_in[`VWidth*(`APPRam_depth*23+74)-1:`VWidth*(`APPRam_depth*23+73)],data_in[`VWidth*(`APPRam_depth*22+74)-1:`VWidth*(`APPRam_depth*22+73)],data_in[`VWidth*(`APPRam_depth*21+74)-1:`VWidth*(`APPRam_depth*21+73)],data_in[`VWidth*(`APPRam_depth*20+74)-1:`VWidth*(`APPRam_depth*20+73)],data_in[`VWidth*(`APPRam_depth*19+74)-1:`VWidth*(`APPRam_depth*19+73)],data_in[`VWidth*(`APPRam_depth*18+74)-1:`VWidth*(`APPRam_depth*18+73)],data_in[`VWidth*(`APPRam_depth*17+74)-1:`VWidth*(`APPRam_depth*17+73)],data_in[`VWidth*(`APPRam_depth*16+74)-1:`VWidth*(`APPRam_depth*16+73)],data_in[`VWidth*(`APPRam_depth*15+74)-1:`VWidth*(`APPRam_depth*15+73)],data_in[`VWidth*(`APPRam_depth*14+74)-1:`VWidth*(`APPRam_depth*14+73)],data_in[`VWidth*(`APPRam_depth*13+74)-1:`VWidth*(`APPRam_depth*13+73)],data_in[`VWidth*(`APPRam_depth*12+74)-1:`VWidth*(`APPRam_depth*12+73)],data_in[`VWidth*(`APPRam_depth*11+74)-1:`VWidth*(`APPRam_depth*11+73)],data_in[`VWidth*(`APPRam_depth*10+74)-1:`VWidth*(`APPRam_depth*10+73)],data_in[`VWidth*(`APPRam_depth*9+74)-1:`VWidth*(`APPRam_depth*9+73)],data_in[`VWidth*(`APPRam_depth*8+74)-1:`VWidth*(`APPRam_depth*8+73)],data_in[`VWidth*(`APPRam_depth*7+74)-1:`VWidth*(`APPRam_depth*7+73)],data_in[`VWidth*(`APPRam_depth*6+74)-1:`VWidth*(`APPRam_depth*6+73)],data_in[`VWidth*(`APPRam_depth*5+74)-1:`VWidth*(`APPRam_depth*5+73)],data_in[`VWidth*(`APPRam_depth*4+74)-1:`VWidth*(`APPRam_depth*4+73)],data_in[`VWidth*(`APPRam_depth*3+74)-1:`VWidth*(`APPRam_depth*3+73)],data_in[`VWidth*(`APPRam_depth*2+74)-1:`VWidth*(`APPRam_depth*2+73)],data_in[`VWidth*(`APPRam_depth*1+74)-1:`VWidth*(`APPRam_depth*1+73)],data_in[`VWidth*(`APPRam_depth*0+74)-1:`VWidth*(`APPRam_depth*0+73)]};
			end
			74:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+75)-1:`VWidth*(`APPRam_depth*31+74)],data_in[`VWidth*(`APPRam_depth*30+75)-1:`VWidth*(`APPRam_depth*30+74)],data_in[`VWidth*(`APPRam_depth*29+75)-1:`VWidth*(`APPRam_depth*29+74)],data_in[`VWidth*(`APPRam_depth*28+75)-1:`VWidth*(`APPRam_depth*28+74)],data_in[`VWidth*(`APPRam_depth*27+75)-1:`VWidth*(`APPRam_depth*27+74)],data_in[`VWidth*(`APPRam_depth*26+75)-1:`VWidth*(`APPRam_depth*26+74)],data_in[`VWidth*(`APPRam_depth*25+75)-1:`VWidth*(`APPRam_depth*25+74)],data_in[`VWidth*(`APPRam_depth*24+75)-1:`VWidth*(`APPRam_depth*24+74)],data_in[`VWidth*(`APPRam_depth*23+75)-1:`VWidth*(`APPRam_depth*23+74)],data_in[`VWidth*(`APPRam_depth*22+75)-1:`VWidth*(`APPRam_depth*22+74)],data_in[`VWidth*(`APPRam_depth*21+75)-1:`VWidth*(`APPRam_depth*21+74)],data_in[`VWidth*(`APPRam_depth*20+75)-1:`VWidth*(`APPRam_depth*20+74)],data_in[`VWidth*(`APPRam_depth*19+75)-1:`VWidth*(`APPRam_depth*19+74)],data_in[`VWidth*(`APPRam_depth*18+75)-1:`VWidth*(`APPRam_depth*18+74)],data_in[`VWidth*(`APPRam_depth*17+75)-1:`VWidth*(`APPRam_depth*17+74)],data_in[`VWidth*(`APPRam_depth*16+75)-1:`VWidth*(`APPRam_depth*16+74)],data_in[`VWidth*(`APPRam_depth*15+75)-1:`VWidth*(`APPRam_depth*15+74)],data_in[`VWidth*(`APPRam_depth*14+75)-1:`VWidth*(`APPRam_depth*14+74)],data_in[`VWidth*(`APPRam_depth*13+75)-1:`VWidth*(`APPRam_depth*13+74)],data_in[`VWidth*(`APPRam_depth*12+75)-1:`VWidth*(`APPRam_depth*12+74)],data_in[`VWidth*(`APPRam_depth*11+75)-1:`VWidth*(`APPRam_depth*11+74)],data_in[`VWidth*(`APPRam_depth*10+75)-1:`VWidth*(`APPRam_depth*10+74)],data_in[`VWidth*(`APPRam_depth*9+75)-1:`VWidth*(`APPRam_depth*9+74)],data_in[`VWidth*(`APPRam_depth*8+75)-1:`VWidth*(`APPRam_depth*8+74)],data_in[`VWidth*(`APPRam_depth*7+75)-1:`VWidth*(`APPRam_depth*7+74)],data_in[`VWidth*(`APPRam_depth*6+75)-1:`VWidth*(`APPRam_depth*6+74)],data_in[`VWidth*(`APPRam_depth*5+75)-1:`VWidth*(`APPRam_depth*5+74)],data_in[`VWidth*(`APPRam_depth*4+75)-1:`VWidth*(`APPRam_depth*4+74)],data_in[`VWidth*(`APPRam_depth*3+75)-1:`VWidth*(`APPRam_depth*3+74)],data_in[`VWidth*(`APPRam_depth*2+75)-1:`VWidth*(`APPRam_depth*2+74)],data_in[`VWidth*(`APPRam_depth*1+75)-1:`VWidth*(`APPRam_depth*1+74)],data_in[`VWidth*(`APPRam_depth*0+75)-1:`VWidth*(`APPRam_depth*0+74)]};
			end
			75:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+76)-1:`VWidth*(`APPRam_depth*31+75)],data_in[`VWidth*(`APPRam_depth*30+76)-1:`VWidth*(`APPRam_depth*30+75)],data_in[`VWidth*(`APPRam_depth*29+76)-1:`VWidth*(`APPRam_depth*29+75)],data_in[`VWidth*(`APPRam_depth*28+76)-1:`VWidth*(`APPRam_depth*28+75)],data_in[`VWidth*(`APPRam_depth*27+76)-1:`VWidth*(`APPRam_depth*27+75)],data_in[`VWidth*(`APPRam_depth*26+76)-1:`VWidth*(`APPRam_depth*26+75)],data_in[`VWidth*(`APPRam_depth*25+76)-1:`VWidth*(`APPRam_depth*25+75)],data_in[`VWidth*(`APPRam_depth*24+76)-1:`VWidth*(`APPRam_depth*24+75)],data_in[`VWidth*(`APPRam_depth*23+76)-1:`VWidth*(`APPRam_depth*23+75)],data_in[`VWidth*(`APPRam_depth*22+76)-1:`VWidth*(`APPRam_depth*22+75)],data_in[`VWidth*(`APPRam_depth*21+76)-1:`VWidth*(`APPRam_depth*21+75)],data_in[`VWidth*(`APPRam_depth*20+76)-1:`VWidth*(`APPRam_depth*20+75)],data_in[`VWidth*(`APPRam_depth*19+76)-1:`VWidth*(`APPRam_depth*19+75)],data_in[`VWidth*(`APPRam_depth*18+76)-1:`VWidth*(`APPRam_depth*18+75)],data_in[`VWidth*(`APPRam_depth*17+76)-1:`VWidth*(`APPRam_depth*17+75)],data_in[`VWidth*(`APPRam_depth*16+76)-1:`VWidth*(`APPRam_depth*16+75)],data_in[`VWidth*(`APPRam_depth*15+76)-1:`VWidth*(`APPRam_depth*15+75)],data_in[`VWidth*(`APPRam_depth*14+76)-1:`VWidth*(`APPRam_depth*14+75)],data_in[`VWidth*(`APPRam_depth*13+76)-1:`VWidth*(`APPRam_depth*13+75)],data_in[`VWidth*(`APPRam_depth*12+76)-1:`VWidth*(`APPRam_depth*12+75)],data_in[`VWidth*(`APPRam_depth*11+76)-1:`VWidth*(`APPRam_depth*11+75)],data_in[`VWidth*(`APPRam_depth*10+76)-1:`VWidth*(`APPRam_depth*10+75)],data_in[`VWidth*(`APPRam_depth*9+76)-1:`VWidth*(`APPRam_depth*9+75)],data_in[`VWidth*(`APPRam_depth*8+76)-1:`VWidth*(`APPRam_depth*8+75)],data_in[`VWidth*(`APPRam_depth*7+76)-1:`VWidth*(`APPRam_depth*7+75)],data_in[`VWidth*(`APPRam_depth*6+76)-1:`VWidth*(`APPRam_depth*6+75)],data_in[`VWidth*(`APPRam_depth*5+76)-1:`VWidth*(`APPRam_depth*5+75)],data_in[`VWidth*(`APPRam_depth*4+76)-1:`VWidth*(`APPRam_depth*4+75)],data_in[`VWidth*(`APPRam_depth*3+76)-1:`VWidth*(`APPRam_depth*3+75)],data_in[`VWidth*(`APPRam_depth*2+76)-1:`VWidth*(`APPRam_depth*2+75)],data_in[`VWidth*(`APPRam_depth*1+76)-1:`VWidth*(`APPRam_depth*1+75)],data_in[`VWidth*(`APPRam_depth*0+76)-1:`VWidth*(`APPRam_depth*0+75)]};
			end
			76:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+77)-1:`VWidth*(`APPRam_depth*31+76)],data_in[`VWidth*(`APPRam_depth*30+77)-1:`VWidth*(`APPRam_depth*30+76)],data_in[`VWidth*(`APPRam_depth*29+77)-1:`VWidth*(`APPRam_depth*29+76)],data_in[`VWidth*(`APPRam_depth*28+77)-1:`VWidth*(`APPRam_depth*28+76)],data_in[`VWidth*(`APPRam_depth*27+77)-1:`VWidth*(`APPRam_depth*27+76)],data_in[`VWidth*(`APPRam_depth*26+77)-1:`VWidth*(`APPRam_depth*26+76)],data_in[`VWidth*(`APPRam_depth*25+77)-1:`VWidth*(`APPRam_depth*25+76)],data_in[`VWidth*(`APPRam_depth*24+77)-1:`VWidth*(`APPRam_depth*24+76)],data_in[`VWidth*(`APPRam_depth*23+77)-1:`VWidth*(`APPRam_depth*23+76)],data_in[`VWidth*(`APPRam_depth*22+77)-1:`VWidth*(`APPRam_depth*22+76)],data_in[`VWidth*(`APPRam_depth*21+77)-1:`VWidth*(`APPRam_depth*21+76)],data_in[`VWidth*(`APPRam_depth*20+77)-1:`VWidth*(`APPRam_depth*20+76)],data_in[`VWidth*(`APPRam_depth*19+77)-1:`VWidth*(`APPRam_depth*19+76)],data_in[`VWidth*(`APPRam_depth*18+77)-1:`VWidth*(`APPRam_depth*18+76)],data_in[`VWidth*(`APPRam_depth*17+77)-1:`VWidth*(`APPRam_depth*17+76)],data_in[`VWidth*(`APPRam_depth*16+77)-1:`VWidth*(`APPRam_depth*16+76)],data_in[`VWidth*(`APPRam_depth*15+77)-1:`VWidth*(`APPRam_depth*15+76)],data_in[`VWidth*(`APPRam_depth*14+77)-1:`VWidth*(`APPRam_depth*14+76)],data_in[`VWidth*(`APPRam_depth*13+77)-1:`VWidth*(`APPRam_depth*13+76)],data_in[`VWidth*(`APPRam_depth*12+77)-1:`VWidth*(`APPRam_depth*12+76)],data_in[`VWidth*(`APPRam_depth*11+77)-1:`VWidth*(`APPRam_depth*11+76)],data_in[`VWidth*(`APPRam_depth*10+77)-1:`VWidth*(`APPRam_depth*10+76)],data_in[`VWidth*(`APPRam_depth*9+77)-1:`VWidth*(`APPRam_depth*9+76)],data_in[`VWidth*(`APPRam_depth*8+77)-1:`VWidth*(`APPRam_depth*8+76)],data_in[`VWidth*(`APPRam_depth*7+77)-1:`VWidth*(`APPRam_depth*7+76)],data_in[`VWidth*(`APPRam_depth*6+77)-1:`VWidth*(`APPRam_depth*6+76)],data_in[`VWidth*(`APPRam_depth*5+77)-1:`VWidth*(`APPRam_depth*5+76)],data_in[`VWidth*(`APPRam_depth*4+77)-1:`VWidth*(`APPRam_depth*4+76)],data_in[`VWidth*(`APPRam_depth*3+77)-1:`VWidth*(`APPRam_depth*3+76)],data_in[`VWidth*(`APPRam_depth*2+77)-1:`VWidth*(`APPRam_depth*2+76)],data_in[`VWidth*(`APPRam_depth*1+77)-1:`VWidth*(`APPRam_depth*1+76)],data_in[`VWidth*(`APPRam_depth*0+77)-1:`VWidth*(`APPRam_depth*0+76)]};
			end
			77:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+78)-1:`VWidth*(`APPRam_depth*31+77)],data_in[`VWidth*(`APPRam_depth*30+78)-1:`VWidth*(`APPRam_depth*30+77)],data_in[`VWidth*(`APPRam_depth*29+78)-1:`VWidth*(`APPRam_depth*29+77)],data_in[`VWidth*(`APPRam_depth*28+78)-1:`VWidth*(`APPRam_depth*28+77)],data_in[`VWidth*(`APPRam_depth*27+78)-1:`VWidth*(`APPRam_depth*27+77)],data_in[`VWidth*(`APPRam_depth*26+78)-1:`VWidth*(`APPRam_depth*26+77)],data_in[`VWidth*(`APPRam_depth*25+78)-1:`VWidth*(`APPRam_depth*25+77)],data_in[`VWidth*(`APPRam_depth*24+78)-1:`VWidth*(`APPRam_depth*24+77)],data_in[`VWidth*(`APPRam_depth*23+78)-1:`VWidth*(`APPRam_depth*23+77)],data_in[`VWidth*(`APPRam_depth*22+78)-1:`VWidth*(`APPRam_depth*22+77)],data_in[`VWidth*(`APPRam_depth*21+78)-1:`VWidth*(`APPRam_depth*21+77)],data_in[`VWidth*(`APPRam_depth*20+78)-1:`VWidth*(`APPRam_depth*20+77)],data_in[`VWidth*(`APPRam_depth*19+78)-1:`VWidth*(`APPRam_depth*19+77)],data_in[`VWidth*(`APPRam_depth*18+78)-1:`VWidth*(`APPRam_depth*18+77)],data_in[`VWidth*(`APPRam_depth*17+78)-1:`VWidth*(`APPRam_depth*17+77)],data_in[`VWidth*(`APPRam_depth*16+78)-1:`VWidth*(`APPRam_depth*16+77)],data_in[`VWidth*(`APPRam_depth*15+78)-1:`VWidth*(`APPRam_depth*15+77)],data_in[`VWidth*(`APPRam_depth*14+78)-1:`VWidth*(`APPRam_depth*14+77)],data_in[`VWidth*(`APPRam_depth*13+78)-1:`VWidth*(`APPRam_depth*13+77)],data_in[`VWidth*(`APPRam_depth*12+78)-1:`VWidth*(`APPRam_depth*12+77)],data_in[`VWidth*(`APPRam_depth*11+78)-1:`VWidth*(`APPRam_depth*11+77)],data_in[`VWidth*(`APPRam_depth*10+78)-1:`VWidth*(`APPRam_depth*10+77)],data_in[`VWidth*(`APPRam_depth*9+78)-1:`VWidth*(`APPRam_depth*9+77)],data_in[`VWidth*(`APPRam_depth*8+78)-1:`VWidth*(`APPRam_depth*8+77)],data_in[`VWidth*(`APPRam_depth*7+78)-1:`VWidth*(`APPRam_depth*7+77)],data_in[`VWidth*(`APPRam_depth*6+78)-1:`VWidth*(`APPRam_depth*6+77)],data_in[`VWidth*(`APPRam_depth*5+78)-1:`VWidth*(`APPRam_depth*5+77)],data_in[`VWidth*(`APPRam_depth*4+78)-1:`VWidth*(`APPRam_depth*4+77)],data_in[`VWidth*(`APPRam_depth*3+78)-1:`VWidth*(`APPRam_depth*3+77)],data_in[`VWidth*(`APPRam_depth*2+78)-1:`VWidth*(`APPRam_depth*2+77)],data_in[`VWidth*(`APPRam_depth*1+78)-1:`VWidth*(`APPRam_depth*1+77)],data_in[`VWidth*(`APPRam_depth*0+78)-1:`VWidth*(`APPRam_depth*0+77)]};
			end
			78:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+79)-1:`VWidth*(`APPRam_depth*31+78)],data_in[`VWidth*(`APPRam_depth*30+79)-1:`VWidth*(`APPRam_depth*30+78)],data_in[`VWidth*(`APPRam_depth*29+79)-1:`VWidth*(`APPRam_depth*29+78)],data_in[`VWidth*(`APPRam_depth*28+79)-1:`VWidth*(`APPRam_depth*28+78)],data_in[`VWidth*(`APPRam_depth*27+79)-1:`VWidth*(`APPRam_depth*27+78)],data_in[`VWidth*(`APPRam_depth*26+79)-1:`VWidth*(`APPRam_depth*26+78)],data_in[`VWidth*(`APPRam_depth*25+79)-1:`VWidth*(`APPRam_depth*25+78)],data_in[`VWidth*(`APPRam_depth*24+79)-1:`VWidth*(`APPRam_depth*24+78)],data_in[`VWidth*(`APPRam_depth*23+79)-1:`VWidth*(`APPRam_depth*23+78)],data_in[`VWidth*(`APPRam_depth*22+79)-1:`VWidth*(`APPRam_depth*22+78)],data_in[`VWidth*(`APPRam_depth*21+79)-1:`VWidth*(`APPRam_depth*21+78)],data_in[`VWidth*(`APPRam_depth*20+79)-1:`VWidth*(`APPRam_depth*20+78)],data_in[`VWidth*(`APPRam_depth*19+79)-1:`VWidth*(`APPRam_depth*19+78)],data_in[`VWidth*(`APPRam_depth*18+79)-1:`VWidth*(`APPRam_depth*18+78)],data_in[`VWidth*(`APPRam_depth*17+79)-1:`VWidth*(`APPRam_depth*17+78)],data_in[`VWidth*(`APPRam_depth*16+79)-1:`VWidth*(`APPRam_depth*16+78)],data_in[`VWidth*(`APPRam_depth*15+79)-1:`VWidth*(`APPRam_depth*15+78)],data_in[`VWidth*(`APPRam_depth*14+79)-1:`VWidth*(`APPRam_depth*14+78)],data_in[`VWidth*(`APPRam_depth*13+79)-1:`VWidth*(`APPRam_depth*13+78)],data_in[`VWidth*(`APPRam_depth*12+79)-1:`VWidth*(`APPRam_depth*12+78)],data_in[`VWidth*(`APPRam_depth*11+79)-1:`VWidth*(`APPRam_depth*11+78)],data_in[`VWidth*(`APPRam_depth*10+79)-1:`VWidth*(`APPRam_depth*10+78)],data_in[`VWidth*(`APPRam_depth*9+79)-1:`VWidth*(`APPRam_depth*9+78)],data_in[`VWidth*(`APPRam_depth*8+79)-1:`VWidth*(`APPRam_depth*8+78)],data_in[`VWidth*(`APPRam_depth*7+79)-1:`VWidth*(`APPRam_depth*7+78)],data_in[`VWidth*(`APPRam_depth*6+79)-1:`VWidth*(`APPRam_depth*6+78)],data_in[`VWidth*(`APPRam_depth*5+79)-1:`VWidth*(`APPRam_depth*5+78)],data_in[`VWidth*(`APPRam_depth*4+79)-1:`VWidth*(`APPRam_depth*4+78)],data_in[`VWidth*(`APPRam_depth*3+79)-1:`VWidth*(`APPRam_depth*3+78)],data_in[`VWidth*(`APPRam_depth*2+79)-1:`VWidth*(`APPRam_depth*2+78)],data_in[`VWidth*(`APPRam_depth*1+79)-1:`VWidth*(`APPRam_depth*1+78)],data_in[`VWidth*(`APPRam_depth*0+79)-1:`VWidth*(`APPRam_depth*0+78)]};
			end
			79:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+80)-1:`VWidth*(`APPRam_depth*31+79)],data_in[`VWidth*(`APPRam_depth*30+80)-1:`VWidth*(`APPRam_depth*30+79)],data_in[`VWidth*(`APPRam_depth*29+80)-1:`VWidth*(`APPRam_depth*29+79)],data_in[`VWidth*(`APPRam_depth*28+80)-1:`VWidth*(`APPRam_depth*28+79)],data_in[`VWidth*(`APPRam_depth*27+80)-1:`VWidth*(`APPRam_depth*27+79)],data_in[`VWidth*(`APPRam_depth*26+80)-1:`VWidth*(`APPRam_depth*26+79)],data_in[`VWidth*(`APPRam_depth*25+80)-1:`VWidth*(`APPRam_depth*25+79)],data_in[`VWidth*(`APPRam_depth*24+80)-1:`VWidth*(`APPRam_depth*24+79)],data_in[`VWidth*(`APPRam_depth*23+80)-1:`VWidth*(`APPRam_depth*23+79)],data_in[`VWidth*(`APPRam_depth*22+80)-1:`VWidth*(`APPRam_depth*22+79)],data_in[`VWidth*(`APPRam_depth*21+80)-1:`VWidth*(`APPRam_depth*21+79)],data_in[`VWidth*(`APPRam_depth*20+80)-1:`VWidth*(`APPRam_depth*20+79)],data_in[`VWidth*(`APPRam_depth*19+80)-1:`VWidth*(`APPRam_depth*19+79)],data_in[`VWidth*(`APPRam_depth*18+80)-1:`VWidth*(`APPRam_depth*18+79)],data_in[`VWidth*(`APPRam_depth*17+80)-1:`VWidth*(`APPRam_depth*17+79)],data_in[`VWidth*(`APPRam_depth*16+80)-1:`VWidth*(`APPRam_depth*16+79)],data_in[`VWidth*(`APPRam_depth*15+80)-1:`VWidth*(`APPRam_depth*15+79)],data_in[`VWidth*(`APPRam_depth*14+80)-1:`VWidth*(`APPRam_depth*14+79)],data_in[`VWidth*(`APPRam_depth*13+80)-1:`VWidth*(`APPRam_depth*13+79)],data_in[`VWidth*(`APPRam_depth*12+80)-1:`VWidth*(`APPRam_depth*12+79)],data_in[`VWidth*(`APPRam_depth*11+80)-1:`VWidth*(`APPRam_depth*11+79)],data_in[`VWidth*(`APPRam_depth*10+80)-1:`VWidth*(`APPRam_depth*10+79)],data_in[`VWidth*(`APPRam_depth*9+80)-1:`VWidth*(`APPRam_depth*9+79)],data_in[`VWidth*(`APPRam_depth*8+80)-1:`VWidth*(`APPRam_depth*8+79)],data_in[`VWidth*(`APPRam_depth*7+80)-1:`VWidth*(`APPRam_depth*7+79)],data_in[`VWidth*(`APPRam_depth*6+80)-1:`VWidth*(`APPRam_depth*6+79)],data_in[`VWidth*(`APPRam_depth*5+80)-1:`VWidth*(`APPRam_depth*5+79)],data_in[`VWidth*(`APPRam_depth*4+80)-1:`VWidth*(`APPRam_depth*4+79)],data_in[`VWidth*(`APPRam_depth*3+80)-1:`VWidth*(`APPRam_depth*3+79)],data_in[`VWidth*(`APPRam_depth*2+80)-1:`VWidth*(`APPRam_depth*2+79)],data_in[`VWidth*(`APPRam_depth*1+80)-1:`VWidth*(`APPRam_depth*1+79)],data_in[`VWidth*(`APPRam_depth*0+80)-1:`VWidth*(`APPRam_depth*0+79)]};
			end
			80:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+81)-1:`VWidth*(`APPRam_depth*31+80)],data_in[`VWidth*(`APPRam_depth*30+81)-1:`VWidth*(`APPRam_depth*30+80)],data_in[`VWidth*(`APPRam_depth*29+81)-1:`VWidth*(`APPRam_depth*29+80)],data_in[`VWidth*(`APPRam_depth*28+81)-1:`VWidth*(`APPRam_depth*28+80)],data_in[`VWidth*(`APPRam_depth*27+81)-1:`VWidth*(`APPRam_depth*27+80)],data_in[`VWidth*(`APPRam_depth*26+81)-1:`VWidth*(`APPRam_depth*26+80)],data_in[`VWidth*(`APPRam_depth*25+81)-1:`VWidth*(`APPRam_depth*25+80)],data_in[`VWidth*(`APPRam_depth*24+81)-1:`VWidth*(`APPRam_depth*24+80)],data_in[`VWidth*(`APPRam_depth*23+81)-1:`VWidth*(`APPRam_depth*23+80)],data_in[`VWidth*(`APPRam_depth*22+81)-1:`VWidth*(`APPRam_depth*22+80)],data_in[`VWidth*(`APPRam_depth*21+81)-1:`VWidth*(`APPRam_depth*21+80)],data_in[`VWidth*(`APPRam_depth*20+81)-1:`VWidth*(`APPRam_depth*20+80)],data_in[`VWidth*(`APPRam_depth*19+81)-1:`VWidth*(`APPRam_depth*19+80)],data_in[`VWidth*(`APPRam_depth*18+81)-1:`VWidth*(`APPRam_depth*18+80)],data_in[`VWidth*(`APPRam_depth*17+81)-1:`VWidth*(`APPRam_depth*17+80)],data_in[`VWidth*(`APPRam_depth*16+81)-1:`VWidth*(`APPRam_depth*16+80)],data_in[`VWidth*(`APPRam_depth*15+81)-1:`VWidth*(`APPRam_depth*15+80)],data_in[`VWidth*(`APPRam_depth*14+81)-1:`VWidth*(`APPRam_depth*14+80)],data_in[`VWidth*(`APPRam_depth*13+81)-1:`VWidth*(`APPRam_depth*13+80)],data_in[`VWidth*(`APPRam_depth*12+81)-1:`VWidth*(`APPRam_depth*12+80)],data_in[`VWidth*(`APPRam_depth*11+81)-1:`VWidth*(`APPRam_depth*11+80)],data_in[`VWidth*(`APPRam_depth*10+81)-1:`VWidth*(`APPRam_depth*10+80)],data_in[`VWidth*(`APPRam_depth*9+81)-1:`VWidth*(`APPRam_depth*9+80)],data_in[`VWidth*(`APPRam_depth*8+81)-1:`VWidth*(`APPRam_depth*8+80)],data_in[`VWidth*(`APPRam_depth*7+81)-1:`VWidth*(`APPRam_depth*7+80)],data_in[`VWidth*(`APPRam_depth*6+81)-1:`VWidth*(`APPRam_depth*6+80)],data_in[`VWidth*(`APPRam_depth*5+81)-1:`VWidth*(`APPRam_depth*5+80)],data_in[`VWidth*(`APPRam_depth*4+81)-1:`VWidth*(`APPRam_depth*4+80)],data_in[`VWidth*(`APPRam_depth*3+81)-1:`VWidth*(`APPRam_depth*3+80)],data_in[`VWidth*(`APPRam_depth*2+81)-1:`VWidth*(`APPRam_depth*2+80)],data_in[`VWidth*(`APPRam_depth*1+81)-1:`VWidth*(`APPRam_depth*1+80)],data_in[`VWidth*(`APPRam_depth*0+81)-1:`VWidth*(`APPRam_depth*0+80)]};
			end
			81:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+82)-1:`VWidth*(`APPRam_depth*31+81)],data_in[`VWidth*(`APPRam_depth*30+82)-1:`VWidth*(`APPRam_depth*30+81)],data_in[`VWidth*(`APPRam_depth*29+82)-1:`VWidth*(`APPRam_depth*29+81)],data_in[`VWidth*(`APPRam_depth*28+82)-1:`VWidth*(`APPRam_depth*28+81)],data_in[`VWidth*(`APPRam_depth*27+82)-1:`VWidth*(`APPRam_depth*27+81)],data_in[`VWidth*(`APPRam_depth*26+82)-1:`VWidth*(`APPRam_depth*26+81)],data_in[`VWidth*(`APPRam_depth*25+82)-1:`VWidth*(`APPRam_depth*25+81)],data_in[`VWidth*(`APPRam_depth*24+82)-1:`VWidth*(`APPRam_depth*24+81)],data_in[`VWidth*(`APPRam_depth*23+82)-1:`VWidth*(`APPRam_depth*23+81)],data_in[`VWidth*(`APPRam_depth*22+82)-1:`VWidth*(`APPRam_depth*22+81)],data_in[`VWidth*(`APPRam_depth*21+82)-1:`VWidth*(`APPRam_depth*21+81)],data_in[`VWidth*(`APPRam_depth*20+82)-1:`VWidth*(`APPRam_depth*20+81)],data_in[`VWidth*(`APPRam_depth*19+82)-1:`VWidth*(`APPRam_depth*19+81)],data_in[`VWidth*(`APPRam_depth*18+82)-1:`VWidth*(`APPRam_depth*18+81)],data_in[`VWidth*(`APPRam_depth*17+82)-1:`VWidth*(`APPRam_depth*17+81)],data_in[`VWidth*(`APPRam_depth*16+82)-1:`VWidth*(`APPRam_depth*16+81)],data_in[`VWidth*(`APPRam_depth*15+82)-1:`VWidth*(`APPRam_depth*15+81)],data_in[`VWidth*(`APPRam_depth*14+82)-1:`VWidth*(`APPRam_depth*14+81)],data_in[`VWidth*(`APPRam_depth*13+82)-1:`VWidth*(`APPRam_depth*13+81)],data_in[`VWidth*(`APPRam_depth*12+82)-1:`VWidth*(`APPRam_depth*12+81)],data_in[`VWidth*(`APPRam_depth*11+82)-1:`VWidth*(`APPRam_depth*11+81)],data_in[`VWidth*(`APPRam_depth*10+82)-1:`VWidth*(`APPRam_depth*10+81)],data_in[`VWidth*(`APPRam_depth*9+82)-1:`VWidth*(`APPRam_depth*9+81)],data_in[`VWidth*(`APPRam_depth*8+82)-1:`VWidth*(`APPRam_depth*8+81)],data_in[`VWidth*(`APPRam_depth*7+82)-1:`VWidth*(`APPRam_depth*7+81)],data_in[`VWidth*(`APPRam_depth*6+82)-1:`VWidth*(`APPRam_depth*6+81)],data_in[`VWidth*(`APPRam_depth*5+82)-1:`VWidth*(`APPRam_depth*5+81)],data_in[`VWidth*(`APPRam_depth*4+82)-1:`VWidth*(`APPRam_depth*4+81)],data_in[`VWidth*(`APPRam_depth*3+82)-1:`VWidth*(`APPRam_depth*3+81)],data_in[`VWidth*(`APPRam_depth*2+82)-1:`VWidth*(`APPRam_depth*2+81)],data_in[`VWidth*(`APPRam_depth*1+82)-1:`VWidth*(`APPRam_depth*1+81)],data_in[`VWidth*(`APPRam_depth*0+82)-1:`VWidth*(`APPRam_depth*0+81)]};
			end
			82:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+83)-1:`VWidth*(`APPRam_depth*31+82)],data_in[`VWidth*(`APPRam_depth*30+83)-1:`VWidth*(`APPRam_depth*30+82)],data_in[`VWidth*(`APPRam_depth*29+83)-1:`VWidth*(`APPRam_depth*29+82)],data_in[`VWidth*(`APPRam_depth*28+83)-1:`VWidth*(`APPRam_depth*28+82)],data_in[`VWidth*(`APPRam_depth*27+83)-1:`VWidth*(`APPRam_depth*27+82)],data_in[`VWidth*(`APPRam_depth*26+83)-1:`VWidth*(`APPRam_depth*26+82)],data_in[`VWidth*(`APPRam_depth*25+83)-1:`VWidth*(`APPRam_depth*25+82)],data_in[`VWidth*(`APPRam_depth*24+83)-1:`VWidth*(`APPRam_depth*24+82)],data_in[`VWidth*(`APPRam_depth*23+83)-1:`VWidth*(`APPRam_depth*23+82)],data_in[`VWidth*(`APPRam_depth*22+83)-1:`VWidth*(`APPRam_depth*22+82)],data_in[`VWidth*(`APPRam_depth*21+83)-1:`VWidth*(`APPRam_depth*21+82)],data_in[`VWidth*(`APPRam_depth*20+83)-1:`VWidth*(`APPRam_depth*20+82)],data_in[`VWidth*(`APPRam_depth*19+83)-1:`VWidth*(`APPRam_depth*19+82)],data_in[`VWidth*(`APPRam_depth*18+83)-1:`VWidth*(`APPRam_depth*18+82)],data_in[`VWidth*(`APPRam_depth*17+83)-1:`VWidth*(`APPRam_depth*17+82)],data_in[`VWidth*(`APPRam_depth*16+83)-1:`VWidth*(`APPRam_depth*16+82)],data_in[`VWidth*(`APPRam_depth*15+83)-1:`VWidth*(`APPRam_depth*15+82)],data_in[`VWidth*(`APPRam_depth*14+83)-1:`VWidth*(`APPRam_depth*14+82)],data_in[`VWidth*(`APPRam_depth*13+83)-1:`VWidth*(`APPRam_depth*13+82)],data_in[`VWidth*(`APPRam_depth*12+83)-1:`VWidth*(`APPRam_depth*12+82)],data_in[`VWidth*(`APPRam_depth*11+83)-1:`VWidth*(`APPRam_depth*11+82)],data_in[`VWidth*(`APPRam_depth*10+83)-1:`VWidth*(`APPRam_depth*10+82)],data_in[`VWidth*(`APPRam_depth*9+83)-1:`VWidth*(`APPRam_depth*9+82)],data_in[`VWidth*(`APPRam_depth*8+83)-1:`VWidth*(`APPRam_depth*8+82)],data_in[`VWidth*(`APPRam_depth*7+83)-1:`VWidth*(`APPRam_depth*7+82)],data_in[`VWidth*(`APPRam_depth*6+83)-1:`VWidth*(`APPRam_depth*6+82)],data_in[`VWidth*(`APPRam_depth*5+83)-1:`VWidth*(`APPRam_depth*5+82)],data_in[`VWidth*(`APPRam_depth*4+83)-1:`VWidth*(`APPRam_depth*4+82)],data_in[`VWidth*(`APPRam_depth*3+83)-1:`VWidth*(`APPRam_depth*3+82)],data_in[`VWidth*(`APPRam_depth*2+83)-1:`VWidth*(`APPRam_depth*2+82)],data_in[`VWidth*(`APPRam_depth*1+83)-1:`VWidth*(`APPRam_depth*1+82)],data_in[`VWidth*(`APPRam_depth*0+83)-1:`VWidth*(`APPRam_depth*0+82)]};
			end
			83:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+84)-1:`VWidth*(`APPRam_depth*31+83)],data_in[`VWidth*(`APPRam_depth*30+84)-1:`VWidth*(`APPRam_depth*30+83)],data_in[`VWidth*(`APPRam_depth*29+84)-1:`VWidth*(`APPRam_depth*29+83)],data_in[`VWidth*(`APPRam_depth*28+84)-1:`VWidth*(`APPRam_depth*28+83)],data_in[`VWidth*(`APPRam_depth*27+84)-1:`VWidth*(`APPRam_depth*27+83)],data_in[`VWidth*(`APPRam_depth*26+84)-1:`VWidth*(`APPRam_depth*26+83)],data_in[`VWidth*(`APPRam_depth*25+84)-1:`VWidth*(`APPRam_depth*25+83)],data_in[`VWidth*(`APPRam_depth*24+84)-1:`VWidth*(`APPRam_depth*24+83)],data_in[`VWidth*(`APPRam_depth*23+84)-1:`VWidth*(`APPRam_depth*23+83)],data_in[`VWidth*(`APPRam_depth*22+84)-1:`VWidth*(`APPRam_depth*22+83)],data_in[`VWidth*(`APPRam_depth*21+84)-1:`VWidth*(`APPRam_depth*21+83)],data_in[`VWidth*(`APPRam_depth*20+84)-1:`VWidth*(`APPRam_depth*20+83)],data_in[`VWidth*(`APPRam_depth*19+84)-1:`VWidth*(`APPRam_depth*19+83)],data_in[`VWidth*(`APPRam_depth*18+84)-1:`VWidth*(`APPRam_depth*18+83)],data_in[`VWidth*(`APPRam_depth*17+84)-1:`VWidth*(`APPRam_depth*17+83)],data_in[`VWidth*(`APPRam_depth*16+84)-1:`VWidth*(`APPRam_depth*16+83)],data_in[`VWidth*(`APPRam_depth*15+84)-1:`VWidth*(`APPRam_depth*15+83)],data_in[`VWidth*(`APPRam_depth*14+84)-1:`VWidth*(`APPRam_depth*14+83)],data_in[`VWidth*(`APPRam_depth*13+84)-1:`VWidth*(`APPRam_depth*13+83)],data_in[`VWidth*(`APPRam_depth*12+84)-1:`VWidth*(`APPRam_depth*12+83)],data_in[`VWidth*(`APPRam_depth*11+84)-1:`VWidth*(`APPRam_depth*11+83)],data_in[`VWidth*(`APPRam_depth*10+84)-1:`VWidth*(`APPRam_depth*10+83)],data_in[`VWidth*(`APPRam_depth*9+84)-1:`VWidth*(`APPRam_depth*9+83)],data_in[`VWidth*(`APPRam_depth*8+84)-1:`VWidth*(`APPRam_depth*8+83)],data_in[`VWidth*(`APPRam_depth*7+84)-1:`VWidth*(`APPRam_depth*7+83)],data_in[`VWidth*(`APPRam_depth*6+84)-1:`VWidth*(`APPRam_depth*6+83)],data_in[`VWidth*(`APPRam_depth*5+84)-1:`VWidth*(`APPRam_depth*5+83)],data_in[`VWidth*(`APPRam_depth*4+84)-1:`VWidth*(`APPRam_depth*4+83)],data_in[`VWidth*(`APPRam_depth*3+84)-1:`VWidth*(`APPRam_depth*3+83)],data_in[`VWidth*(`APPRam_depth*2+84)-1:`VWidth*(`APPRam_depth*2+83)],data_in[`VWidth*(`APPRam_depth*1+84)-1:`VWidth*(`APPRam_depth*1+83)],data_in[`VWidth*(`APPRam_depth*0+84)-1:`VWidth*(`APPRam_depth*0+83)]};
			end
			84:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+85)-1:`VWidth*(`APPRam_depth*31+84)],data_in[`VWidth*(`APPRam_depth*30+85)-1:`VWidth*(`APPRam_depth*30+84)],data_in[`VWidth*(`APPRam_depth*29+85)-1:`VWidth*(`APPRam_depth*29+84)],data_in[`VWidth*(`APPRam_depth*28+85)-1:`VWidth*(`APPRam_depth*28+84)],data_in[`VWidth*(`APPRam_depth*27+85)-1:`VWidth*(`APPRam_depth*27+84)],data_in[`VWidth*(`APPRam_depth*26+85)-1:`VWidth*(`APPRam_depth*26+84)],data_in[`VWidth*(`APPRam_depth*25+85)-1:`VWidth*(`APPRam_depth*25+84)],data_in[`VWidth*(`APPRam_depth*24+85)-1:`VWidth*(`APPRam_depth*24+84)],data_in[`VWidth*(`APPRam_depth*23+85)-1:`VWidth*(`APPRam_depth*23+84)],data_in[`VWidth*(`APPRam_depth*22+85)-1:`VWidth*(`APPRam_depth*22+84)],data_in[`VWidth*(`APPRam_depth*21+85)-1:`VWidth*(`APPRam_depth*21+84)],data_in[`VWidth*(`APPRam_depth*20+85)-1:`VWidth*(`APPRam_depth*20+84)],data_in[`VWidth*(`APPRam_depth*19+85)-1:`VWidth*(`APPRam_depth*19+84)],data_in[`VWidth*(`APPRam_depth*18+85)-1:`VWidth*(`APPRam_depth*18+84)],data_in[`VWidth*(`APPRam_depth*17+85)-1:`VWidth*(`APPRam_depth*17+84)],data_in[`VWidth*(`APPRam_depth*16+85)-1:`VWidth*(`APPRam_depth*16+84)],data_in[`VWidth*(`APPRam_depth*15+85)-1:`VWidth*(`APPRam_depth*15+84)],data_in[`VWidth*(`APPRam_depth*14+85)-1:`VWidth*(`APPRam_depth*14+84)],data_in[`VWidth*(`APPRam_depth*13+85)-1:`VWidth*(`APPRam_depth*13+84)],data_in[`VWidth*(`APPRam_depth*12+85)-1:`VWidth*(`APPRam_depth*12+84)],data_in[`VWidth*(`APPRam_depth*11+85)-1:`VWidth*(`APPRam_depth*11+84)],data_in[`VWidth*(`APPRam_depth*10+85)-1:`VWidth*(`APPRam_depth*10+84)],data_in[`VWidth*(`APPRam_depth*9+85)-1:`VWidth*(`APPRam_depth*9+84)],data_in[`VWidth*(`APPRam_depth*8+85)-1:`VWidth*(`APPRam_depth*8+84)],data_in[`VWidth*(`APPRam_depth*7+85)-1:`VWidth*(`APPRam_depth*7+84)],data_in[`VWidth*(`APPRam_depth*6+85)-1:`VWidth*(`APPRam_depth*6+84)],data_in[`VWidth*(`APPRam_depth*5+85)-1:`VWidth*(`APPRam_depth*5+84)],data_in[`VWidth*(`APPRam_depth*4+85)-1:`VWidth*(`APPRam_depth*4+84)],data_in[`VWidth*(`APPRam_depth*3+85)-1:`VWidth*(`APPRam_depth*3+84)],data_in[`VWidth*(`APPRam_depth*2+85)-1:`VWidth*(`APPRam_depth*2+84)],data_in[`VWidth*(`APPRam_depth*1+85)-1:`VWidth*(`APPRam_depth*1+84)],data_in[`VWidth*(`APPRam_depth*0+85)-1:`VWidth*(`APPRam_depth*0+84)]};
			end
			85:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+86)-1:`VWidth*(`APPRam_depth*31+85)],data_in[`VWidth*(`APPRam_depth*30+86)-1:`VWidth*(`APPRam_depth*30+85)],data_in[`VWidth*(`APPRam_depth*29+86)-1:`VWidth*(`APPRam_depth*29+85)],data_in[`VWidth*(`APPRam_depth*28+86)-1:`VWidth*(`APPRam_depth*28+85)],data_in[`VWidth*(`APPRam_depth*27+86)-1:`VWidth*(`APPRam_depth*27+85)],data_in[`VWidth*(`APPRam_depth*26+86)-1:`VWidth*(`APPRam_depth*26+85)],data_in[`VWidth*(`APPRam_depth*25+86)-1:`VWidth*(`APPRam_depth*25+85)],data_in[`VWidth*(`APPRam_depth*24+86)-1:`VWidth*(`APPRam_depth*24+85)],data_in[`VWidth*(`APPRam_depth*23+86)-1:`VWidth*(`APPRam_depth*23+85)],data_in[`VWidth*(`APPRam_depth*22+86)-1:`VWidth*(`APPRam_depth*22+85)],data_in[`VWidth*(`APPRam_depth*21+86)-1:`VWidth*(`APPRam_depth*21+85)],data_in[`VWidth*(`APPRam_depth*20+86)-1:`VWidth*(`APPRam_depth*20+85)],data_in[`VWidth*(`APPRam_depth*19+86)-1:`VWidth*(`APPRam_depth*19+85)],data_in[`VWidth*(`APPRam_depth*18+86)-1:`VWidth*(`APPRam_depth*18+85)],data_in[`VWidth*(`APPRam_depth*17+86)-1:`VWidth*(`APPRam_depth*17+85)],data_in[`VWidth*(`APPRam_depth*16+86)-1:`VWidth*(`APPRam_depth*16+85)],data_in[`VWidth*(`APPRam_depth*15+86)-1:`VWidth*(`APPRam_depth*15+85)],data_in[`VWidth*(`APPRam_depth*14+86)-1:`VWidth*(`APPRam_depth*14+85)],data_in[`VWidth*(`APPRam_depth*13+86)-1:`VWidth*(`APPRam_depth*13+85)],data_in[`VWidth*(`APPRam_depth*12+86)-1:`VWidth*(`APPRam_depth*12+85)],data_in[`VWidth*(`APPRam_depth*11+86)-1:`VWidth*(`APPRam_depth*11+85)],data_in[`VWidth*(`APPRam_depth*10+86)-1:`VWidth*(`APPRam_depth*10+85)],data_in[`VWidth*(`APPRam_depth*9+86)-1:`VWidth*(`APPRam_depth*9+85)],data_in[`VWidth*(`APPRam_depth*8+86)-1:`VWidth*(`APPRam_depth*8+85)],data_in[`VWidth*(`APPRam_depth*7+86)-1:`VWidth*(`APPRam_depth*7+85)],data_in[`VWidth*(`APPRam_depth*6+86)-1:`VWidth*(`APPRam_depth*6+85)],data_in[`VWidth*(`APPRam_depth*5+86)-1:`VWidth*(`APPRam_depth*5+85)],data_in[`VWidth*(`APPRam_depth*4+86)-1:`VWidth*(`APPRam_depth*4+85)],data_in[`VWidth*(`APPRam_depth*3+86)-1:`VWidth*(`APPRam_depth*3+85)],data_in[`VWidth*(`APPRam_depth*2+86)-1:`VWidth*(`APPRam_depth*2+85)],data_in[`VWidth*(`APPRam_depth*1+86)-1:`VWidth*(`APPRam_depth*1+85)],data_in[`VWidth*(`APPRam_depth*0+86)-1:`VWidth*(`APPRam_depth*0+85)]};
			end
			86:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+87)-1:`VWidth*(`APPRam_depth*31+86)],data_in[`VWidth*(`APPRam_depth*30+87)-1:`VWidth*(`APPRam_depth*30+86)],data_in[`VWidth*(`APPRam_depth*29+87)-1:`VWidth*(`APPRam_depth*29+86)],data_in[`VWidth*(`APPRam_depth*28+87)-1:`VWidth*(`APPRam_depth*28+86)],data_in[`VWidth*(`APPRam_depth*27+87)-1:`VWidth*(`APPRam_depth*27+86)],data_in[`VWidth*(`APPRam_depth*26+87)-1:`VWidth*(`APPRam_depth*26+86)],data_in[`VWidth*(`APPRam_depth*25+87)-1:`VWidth*(`APPRam_depth*25+86)],data_in[`VWidth*(`APPRam_depth*24+87)-1:`VWidth*(`APPRam_depth*24+86)],data_in[`VWidth*(`APPRam_depth*23+87)-1:`VWidth*(`APPRam_depth*23+86)],data_in[`VWidth*(`APPRam_depth*22+87)-1:`VWidth*(`APPRam_depth*22+86)],data_in[`VWidth*(`APPRam_depth*21+87)-1:`VWidth*(`APPRam_depth*21+86)],data_in[`VWidth*(`APPRam_depth*20+87)-1:`VWidth*(`APPRam_depth*20+86)],data_in[`VWidth*(`APPRam_depth*19+87)-1:`VWidth*(`APPRam_depth*19+86)],data_in[`VWidth*(`APPRam_depth*18+87)-1:`VWidth*(`APPRam_depth*18+86)],data_in[`VWidth*(`APPRam_depth*17+87)-1:`VWidth*(`APPRam_depth*17+86)],data_in[`VWidth*(`APPRam_depth*16+87)-1:`VWidth*(`APPRam_depth*16+86)],data_in[`VWidth*(`APPRam_depth*15+87)-1:`VWidth*(`APPRam_depth*15+86)],data_in[`VWidth*(`APPRam_depth*14+87)-1:`VWidth*(`APPRam_depth*14+86)],data_in[`VWidth*(`APPRam_depth*13+87)-1:`VWidth*(`APPRam_depth*13+86)],data_in[`VWidth*(`APPRam_depth*12+87)-1:`VWidth*(`APPRam_depth*12+86)],data_in[`VWidth*(`APPRam_depth*11+87)-1:`VWidth*(`APPRam_depth*11+86)],data_in[`VWidth*(`APPRam_depth*10+87)-1:`VWidth*(`APPRam_depth*10+86)],data_in[`VWidth*(`APPRam_depth*9+87)-1:`VWidth*(`APPRam_depth*9+86)],data_in[`VWidth*(`APPRam_depth*8+87)-1:`VWidth*(`APPRam_depth*8+86)],data_in[`VWidth*(`APPRam_depth*7+87)-1:`VWidth*(`APPRam_depth*7+86)],data_in[`VWidth*(`APPRam_depth*6+87)-1:`VWidth*(`APPRam_depth*6+86)],data_in[`VWidth*(`APPRam_depth*5+87)-1:`VWidth*(`APPRam_depth*5+86)],data_in[`VWidth*(`APPRam_depth*4+87)-1:`VWidth*(`APPRam_depth*4+86)],data_in[`VWidth*(`APPRam_depth*3+87)-1:`VWidth*(`APPRam_depth*3+86)],data_in[`VWidth*(`APPRam_depth*2+87)-1:`VWidth*(`APPRam_depth*2+86)],data_in[`VWidth*(`APPRam_depth*1+87)-1:`VWidth*(`APPRam_depth*1+86)],data_in[`VWidth*(`APPRam_depth*0+87)-1:`VWidth*(`APPRam_depth*0+86)]};
			end
			87:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+88)-1:`VWidth*(`APPRam_depth*31+87)],data_in[`VWidth*(`APPRam_depth*30+88)-1:`VWidth*(`APPRam_depth*30+87)],data_in[`VWidth*(`APPRam_depth*29+88)-1:`VWidth*(`APPRam_depth*29+87)],data_in[`VWidth*(`APPRam_depth*28+88)-1:`VWidth*(`APPRam_depth*28+87)],data_in[`VWidth*(`APPRam_depth*27+88)-1:`VWidth*(`APPRam_depth*27+87)],data_in[`VWidth*(`APPRam_depth*26+88)-1:`VWidth*(`APPRam_depth*26+87)],data_in[`VWidth*(`APPRam_depth*25+88)-1:`VWidth*(`APPRam_depth*25+87)],data_in[`VWidth*(`APPRam_depth*24+88)-1:`VWidth*(`APPRam_depth*24+87)],data_in[`VWidth*(`APPRam_depth*23+88)-1:`VWidth*(`APPRam_depth*23+87)],data_in[`VWidth*(`APPRam_depth*22+88)-1:`VWidth*(`APPRam_depth*22+87)],data_in[`VWidth*(`APPRam_depth*21+88)-1:`VWidth*(`APPRam_depth*21+87)],data_in[`VWidth*(`APPRam_depth*20+88)-1:`VWidth*(`APPRam_depth*20+87)],data_in[`VWidth*(`APPRam_depth*19+88)-1:`VWidth*(`APPRam_depth*19+87)],data_in[`VWidth*(`APPRam_depth*18+88)-1:`VWidth*(`APPRam_depth*18+87)],data_in[`VWidth*(`APPRam_depth*17+88)-1:`VWidth*(`APPRam_depth*17+87)],data_in[`VWidth*(`APPRam_depth*16+88)-1:`VWidth*(`APPRam_depth*16+87)],data_in[`VWidth*(`APPRam_depth*15+88)-1:`VWidth*(`APPRam_depth*15+87)],data_in[`VWidth*(`APPRam_depth*14+88)-1:`VWidth*(`APPRam_depth*14+87)],data_in[`VWidth*(`APPRam_depth*13+88)-1:`VWidth*(`APPRam_depth*13+87)],data_in[`VWidth*(`APPRam_depth*12+88)-1:`VWidth*(`APPRam_depth*12+87)],data_in[`VWidth*(`APPRam_depth*11+88)-1:`VWidth*(`APPRam_depth*11+87)],data_in[`VWidth*(`APPRam_depth*10+88)-1:`VWidth*(`APPRam_depth*10+87)],data_in[`VWidth*(`APPRam_depth*9+88)-1:`VWidth*(`APPRam_depth*9+87)],data_in[`VWidth*(`APPRam_depth*8+88)-1:`VWidth*(`APPRam_depth*8+87)],data_in[`VWidth*(`APPRam_depth*7+88)-1:`VWidth*(`APPRam_depth*7+87)],data_in[`VWidth*(`APPRam_depth*6+88)-1:`VWidth*(`APPRam_depth*6+87)],data_in[`VWidth*(`APPRam_depth*5+88)-1:`VWidth*(`APPRam_depth*5+87)],data_in[`VWidth*(`APPRam_depth*4+88)-1:`VWidth*(`APPRam_depth*4+87)],data_in[`VWidth*(`APPRam_depth*3+88)-1:`VWidth*(`APPRam_depth*3+87)],data_in[`VWidth*(`APPRam_depth*2+88)-1:`VWidth*(`APPRam_depth*2+87)],data_in[`VWidth*(`APPRam_depth*1+88)-1:`VWidth*(`APPRam_depth*1+87)],data_in[`VWidth*(`APPRam_depth*0+88)-1:`VWidth*(`APPRam_depth*0+87)]};
			end
			88:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+89)-1:`VWidth*(`APPRam_depth*31+88)],data_in[`VWidth*(`APPRam_depth*30+89)-1:`VWidth*(`APPRam_depth*30+88)],data_in[`VWidth*(`APPRam_depth*29+89)-1:`VWidth*(`APPRam_depth*29+88)],data_in[`VWidth*(`APPRam_depth*28+89)-1:`VWidth*(`APPRam_depth*28+88)],data_in[`VWidth*(`APPRam_depth*27+89)-1:`VWidth*(`APPRam_depth*27+88)],data_in[`VWidth*(`APPRam_depth*26+89)-1:`VWidth*(`APPRam_depth*26+88)],data_in[`VWidth*(`APPRam_depth*25+89)-1:`VWidth*(`APPRam_depth*25+88)],data_in[`VWidth*(`APPRam_depth*24+89)-1:`VWidth*(`APPRam_depth*24+88)],data_in[`VWidth*(`APPRam_depth*23+89)-1:`VWidth*(`APPRam_depth*23+88)],data_in[`VWidth*(`APPRam_depth*22+89)-1:`VWidth*(`APPRam_depth*22+88)],data_in[`VWidth*(`APPRam_depth*21+89)-1:`VWidth*(`APPRam_depth*21+88)],data_in[`VWidth*(`APPRam_depth*20+89)-1:`VWidth*(`APPRam_depth*20+88)],data_in[`VWidth*(`APPRam_depth*19+89)-1:`VWidth*(`APPRam_depth*19+88)],data_in[`VWidth*(`APPRam_depth*18+89)-1:`VWidth*(`APPRam_depth*18+88)],data_in[`VWidth*(`APPRam_depth*17+89)-1:`VWidth*(`APPRam_depth*17+88)],data_in[`VWidth*(`APPRam_depth*16+89)-1:`VWidth*(`APPRam_depth*16+88)],data_in[`VWidth*(`APPRam_depth*15+89)-1:`VWidth*(`APPRam_depth*15+88)],data_in[`VWidth*(`APPRam_depth*14+89)-1:`VWidth*(`APPRam_depth*14+88)],data_in[`VWidth*(`APPRam_depth*13+89)-1:`VWidth*(`APPRam_depth*13+88)],data_in[`VWidth*(`APPRam_depth*12+89)-1:`VWidth*(`APPRam_depth*12+88)],data_in[`VWidth*(`APPRam_depth*11+89)-1:`VWidth*(`APPRam_depth*11+88)],data_in[`VWidth*(`APPRam_depth*10+89)-1:`VWidth*(`APPRam_depth*10+88)],data_in[`VWidth*(`APPRam_depth*9+89)-1:`VWidth*(`APPRam_depth*9+88)],data_in[`VWidth*(`APPRam_depth*8+89)-1:`VWidth*(`APPRam_depth*8+88)],data_in[`VWidth*(`APPRam_depth*7+89)-1:`VWidth*(`APPRam_depth*7+88)],data_in[`VWidth*(`APPRam_depth*6+89)-1:`VWidth*(`APPRam_depth*6+88)],data_in[`VWidth*(`APPRam_depth*5+89)-1:`VWidth*(`APPRam_depth*5+88)],data_in[`VWidth*(`APPRam_depth*4+89)-1:`VWidth*(`APPRam_depth*4+88)],data_in[`VWidth*(`APPRam_depth*3+89)-1:`VWidth*(`APPRam_depth*3+88)],data_in[`VWidth*(`APPRam_depth*2+89)-1:`VWidth*(`APPRam_depth*2+88)],data_in[`VWidth*(`APPRam_depth*1+89)-1:`VWidth*(`APPRam_depth*1+88)],data_in[`VWidth*(`APPRam_depth*0+89)-1:`VWidth*(`APPRam_depth*0+88)]};
			end
			89:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+90)-1:`VWidth*(`APPRam_depth*31+89)],data_in[`VWidth*(`APPRam_depth*30+90)-1:`VWidth*(`APPRam_depth*30+89)],data_in[`VWidth*(`APPRam_depth*29+90)-1:`VWidth*(`APPRam_depth*29+89)],data_in[`VWidth*(`APPRam_depth*28+90)-1:`VWidth*(`APPRam_depth*28+89)],data_in[`VWidth*(`APPRam_depth*27+90)-1:`VWidth*(`APPRam_depth*27+89)],data_in[`VWidth*(`APPRam_depth*26+90)-1:`VWidth*(`APPRam_depth*26+89)],data_in[`VWidth*(`APPRam_depth*25+90)-1:`VWidth*(`APPRam_depth*25+89)],data_in[`VWidth*(`APPRam_depth*24+90)-1:`VWidth*(`APPRam_depth*24+89)],data_in[`VWidth*(`APPRam_depth*23+90)-1:`VWidth*(`APPRam_depth*23+89)],data_in[`VWidth*(`APPRam_depth*22+90)-1:`VWidth*(`APPRam_depth*22+89)],data_in[`VWidth*(`APPRam_depth*21+90)-1:`VWidth*(`APPRam_depth*21+89)],data_in[`VWidth*(`APPRam_depth*20+90)-1:`VWidth*(`APPRam_depth*20+89)],data_in[`VWidth*(`APPRam_depth*19+90)-1:`VWidth*(`APPRam_depth*19+89)],data_in[`VWidth*(`APPRam_depth*18+90)-1:`VWidth*(`APPRam_depth*18+89)],data_in[`VWidth*(`APPRam_depth*17+90)-1:`VWidth*(`APPRam_depth*17+89)],data_in[`VWidth*(`APPRam_depth*16+90)-1:`VWidth*(`APPRam_depth*16+89)],data_in[`VWidth*(`APPRam_depth*15+90)-1:`VWidth*(`APPRam_depth*15+89)],data_in[`VWidth*(`APPRam_depth*14+90)-1:`VWidth*(`APPRam_depth*14+89)],data_in[`VWidth*(`APPRam_depth*13+90)-1:`VWidth*(`APPRam_depth*13+89)],data_in[`VWidth*(`APPRam_depth*12+90)-1:`VWidth*(`APPRam_depth*12+89)],data_in[`VWidth*(`APPRam_depth*11+90)-1:`VWidth*(`APPRam_depth*11+89)],data_in[`VWidth*(`APPRam_depth*10+90)-1:`VWidth*(`APPRam_depth*10+89)],data_in[`VWidth*(`APPRam_depth*9+90)-1:`VWidth*(`APPRam_depth*9+89)],data_in[`VWidth*(`APPRam_depth*8+90)-1:`VWidth*(`APPRam_depth*8+89)],data_in[`VWidth*(`APPRam_depth*7+90)-1:`VWidth*(`APPRam_depth*7+89)],data_in[`VWidth*(`APPRam_depth*6+90)-1:`VWidth*(`APPRam_depth*6+89)],data_in[`VWidth*(`APPRam_depth*5+90)-1:`VWidth*(`APPRam_depth*5+89)],data_in[`VWidth*(`APPRam_depth*4+90)-1:`VWidth*(`APPRam_depth*4+89)],data_in[`VWidth*(`APPRam_depth*3+90)-1:`VWidth*(`APPRam_depth*3+89)],data_in[`VWidth*(`APPRam_depth*2+90)-1:`VWidth*(`APPRam_depth*2+89)],data_in[`VWidth*(`APPRam_depth*1+90)-1:`VWidth*(`APPRam_depth*1+89)],data_in[`VWidth*(`APPRam_depth*0+90)-1:`VWidth*(`APPRam_depth*0+89)]};
			end
			90:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+91)-1:`VWidth*(`APPRam_depth*31+90)],data_in[`VWidth*(`APPRam_depth*30+91)-1:`VWidth*(`APPRam_depth*30+90)],data_in[`VWidth*(`APPRam_depth*29+91)-1:`VWidth*(`APPRam_depth*29+90)],data_in[`VWidth*(`APPRam_depth*28+91)-1:`VWidth*(`APPRam_depth*28+90)],data_in[`VWidth*(`APPRam_depth*27+91)-1:`VWidth*(`APPRam_depth*27+90)],data_in[`VWidth*(`APPRam_depth*26+91)-1:`VWidth*(`APPRam_depth*26+90)],data_in[`VWidth*(`APPRam_depth*25+91)-1:`VWidth*(`APPRam_depth*25+90)],data_in[`VWidth*(`APPRam_depth*24+91)-1:`VWidth*(`APPRam_depth*24+90)],data_in[`VWidth*(`APPRam_depth*23+91)-1:`VWidth*(`APPRam_depth*23+90)],data_in[`VWidth*(`APPRam_depth*22+91)-1:`VWidth*(`APPRam_depth*22+90)],data_in[`VWidth*(`APPRam_depth*21+91)-1:`VWidth*(`APPRam_depth*21+90)],data_in[`VWidth*(`APPRam_depth*20+91)-1:`VWidth*(`APPRam_depth*20+90)],data_in[`VWidth*(`APPRam_depth*19+91)-1:`VWidth*(`APPRam_depth*19+90)],data_in[`VWidth*(`APPRam_depth*18+91)-1:`VWidth*(`APPRam_depth*18+90)],data_in[`VWidth*(`APPRam_depth*17+91)-1:`VWidth*(`APPRam_depth*17+90)],data_in[`VWidth*(`APPRam_depth*16+91)-1:`VWidth*(`APPRam_depth*16+90)],data_in[`VWidth*(`APPRam_depth*15+91)-1:`VWidth*(`APPRam_depth*15+90)],data_in[`VWidth*(`APPRam_depth*14+91)-1:`VWidth*(`APPRam_depth*14+90)],data_in[`VWidth*(`APPRam_depth*13+91)-1:`VWidth*(`APPRam_depth*13+90)],data_in[`VWidth*(`APPRam_depth*12+91)-1:`VWidth*(`APPRam_depth*12+90)],data_in[`VWidth*(`APPRam_depth*11+91)-1:`VWidth*(`APPRam_depth*11+90)],data_in[`VWidth*(`APPRam_depth*10+91)-1:`VWidth*(`APPRam_depth*10+90)],data_in[`VWidth*(`APPRam_depth*9+91)-1:`VWidth*(`APPRam_depth*9+90)],data_in[`VWidth*(`APPRam_depth*8+91)-1:`VWidth*(`APPRam_depth*8+90)],data_in[`VWidth*(`APPRam_depth*7+91)-1:`VWidth*(`APPRam_depth*7+90)],data_in[`VWidth*(`APPRam_depth*6+91)-1:`VWidth*(`APPRam_depth*6+90)],data_in[`VWidth*(`APPRam_depth*5+91)-1:`VWidth*(`APPRam_depth*5+90)],data_in[`VWidth*(`APPRam_depth*4+91)-1:`VWidth*(`APPRam_depth*4+90)],data_in[`VWidth*(`APPRam_depth*3+91)-1:`VWidth*(`APPRam_depth*3+90)],data_in[`VWidth*(`APPRam_depth*2+91)-1:`VWidth*(`APPRam_depth*2+90)],data_in[`VWidth*(`APPRam_depth*1+91)-1:`VWidth*(`APPRam_depth*1+90)],data_in[`VWidth*(`APPRam_depth*0+91)-1:`VWidth*(`APPRam_depth*0+90)]};
			end
			91:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+92)-1:`VWidth*(`APPRam_depth*31+91)],data_in[`VWidth*(`APPRam_depth*30+92)-1:`VWidth*(`APPRam_depth*30+91)],data_in[`VWidth*(`APPRam_depth*29+92)-1:`VWidth*(`APPRam_depth*29+91)],data_in[`VWidth*(`APPRam_depth*28+92)-1:`VWidth*(`APPRam_depth*28+91)],data_in[`VWidth*(`APPRam_depth*27+92)-1:`VWidth*(`APPRam_depth*27+91)],data_in[`VWidth*(`APPRam_depth*26+92)-1:`VWidth*(`APPRam_depth*26+91)],data_in[`VWidth*(`APPRam_depth*25+92)-1:`VWidth*(`APPRam_depth*25+91)],data_in[`VWidth*(`APPRam_depth*24+92)-1:`VWidth*(`APPRam_depth*24+91)],data_in[`VWidth*(`APPRam_depth*23+92)-1:`VWidth*(`APPRam_depth*23+91)],data_in[`VWidth*(`APPRam_depth*22+92)-1:`VWidth*(`APPRam_depth*22+91)],data_in[`VWidth*(`APPRam_depth*21+92)-1:`VWidth*(`APPRam_depth*21+91)],data_in[`VWidth*(`APPRam_depth*20+92)-1:`VWidth*(`APPRam_depth*20+91)],data_in[`VWidth*(`APPRam_depth*19+92)-1:`VWidth*(`APPRam_depth*19+91)],data_in[`VWidth*(`APPRam_depth*18+92)-1:`VWidth*(`APPRam_depth*18+91)],data_in[`VWidth*(`APPRam_depth*17+92)-1:`VWidth*(`APPRam_depth*17+91)],data_in[`VWidth*(`APPRam_depth*16+92)-1:`VWidth*(`APPRam_depth*16+91)],data_in[`VWidth*(`APPRam_depth*15+92)-1:`VWidth*(`APPRam_depth*15+91)],data_in[`VWidth*(`APPRam_depth*14+92)-1:`VWidth*(`APPRam_depth*14+91)],data_in[`VWidth*(`APPRam_depth*13+92)-1:`VWidth*(`APPRam_depth*13+91)],data_in[`VWidth*(`APPRam_depth*12+92)-1:`VWidth*(`APPRam_depth*12+91)],data_in[`VWidth*(`APPRam_depth*11+92)-1:`VWidth*(`APPRam_depth*11+91)],data_in[`VWidth*(`APPRam_depth*10+92)-1:`VWidth*(`APPRam_depth*10+91)],data_in[`VWidth*(`APPRam_depth*9+92)-1:`VWidth*(`APPRam_depth*9+91)],data_in[`VWidth*(`APPRam_depth*8+92)-1:`VWidth*(`APPRam_depth*8+91)],data_in[`VWidth*(`APPRam_depth*7+92)-1:`VWidth*(`APPRam_depth*7+91)],data_in[`VWidth*(`APPRam_depth*6+92)-1:`VWidth*(`APPRam_depth*6+91)],data_in[`VWidth*(`APPRam_depth*5+92)-1:`VWidth*(`APPRam_depth*5+91)],data_in[`VWidth*(`APPRam_depth*4+92)-1:`VWidth*(`APPRam_depth*4+91)],data_in[`VWidth*(`APPRam_depth*3+92)-1:`VWidth*(`APPRam_depth*3+91)],data_in[`VWidth*(`APPRam_depth*2+92)-1:`VWidth*(`APPRam_depth*2+91)],data_in[`VWidth*(`APPRam_depth*1+92)-1:`VWidth*(`APPRam_depth*1+91)],data_in[`VWidth*(`APPRam_depth*0+92)-1:`VWidth*(`APPRam_depth*0+91)]};
			end
			92:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+93)-1:`VWidth*(`APPRam_depth*31+92)],data_in[`VWidth*(`APPRam_depth*30+93)-1:`VWidth*(`APPRam_depth*30+92)],data_in[`VWidth*(`APPRam_depth*29+93)-1:`VWidth*(`APPRam_depth*29+92)],data_in[`VWidth*(`APPRam_depth*28+93)-1:`VWidth*(`APPRam_depth*28+92)],data_in[`VWidth*(`APPRam_depth*27+93)-1:`VWidth*(`APPRam_depth*27+92)],data_in[`VWidth*(`APPRam_depth*26+93)-1:`VWidth*(`APPRam_depth*26+92)],data_in[`VWidth*(`APPRam_depth*25+93)-1:`VWidth*(`APPRam_depth*25+92)],data_in[`VWidth*(`APPRam_depth*24+93)-1:`VWidth*(`APPRam_depth*24+92)],data_in[`VWidth*(`APPRam_depth*23+93)-1:`VWidth*(`APPRam_depth*23+92)],data_in[`VWidth*(`APPRam_depth*22+93)-1:`VWidth*(`APPRam_depth*22+92)],data_in[`VWidth*(`APPRam_depth*21+93)-1:`VWidth*(`APPRam_depth*21+92)],data_in[`VWidth*(`APPRam_depth*20+93)-1:`VWidth*(`APPRam_depth*20+92)],data_in[`VWidth*(`APPRam_depth*19+93)-1:`VWidth*(`APPRam_depth*19+92)],data_in[`VWidth*(`APPRam_depth*18+93)-1:`VWidth*(`APPRam_depth*18+92)],data_in[`VWidth*(`APPRam_depth*17+93)-1:`VWidth*(`APPRam_depth*17+92)],data_in[`VWidth*(`APPRam_depth*16+93)-1:`VWidth*(`APPRam_depth*16+92)],data_in[`VWidth*(`APPRam_depth*15+93)-1:`VWidth*(`APPRam_depth*15+92)],data_in[`VWidth*(`APPRam_depth*14+93)-1:`VWidth*(`APPRam_depth*14+92)],data_in[`VWidth*(`APPRam_depth*13+93)-1:`VWidth*(`APPRam_depth*13+92)],data_in[`VWidth*(`APPRam_depth*12+93)-1:`VWidth*(`APPRam_depth*12+92)],data_in[`VWidth*(`APPRam_depth*11+93)-1:`VWidth*(`APPRam_depth*11+92)],data_in[`VWidth*(`APPRam_depth*10+93)-1:`VWidth*(`APPRam_depth*10+92)],data_in[`VWidth*(`APPRam_depth*9+93)-1:`VWidth*(`APPRam_depth*9+92)],data_in[`VWidth*(`APPRam_depth*8+93)-1:`VWidth*(`APPRam_depth*8+92)],data_in[`VWidth*(`APPRam_depth*7+93)-1:`VWidth*(`APPRam_depth*7+92)],data_in[`VWidth*(`APPRam_depth*6+93)-1:`VWidth*(`APPRam_depth*6+92)],data_in[`VWidth*(`APPRam_depth*5+93)-1:`VWidth*(`APPRam_depth*5+92)],data_in[`VWidth*(`APPRam_depth*4+93)-1:`VWidth*(`APPRam_depth*4+92)],data_in[`VWidth*(`APPRam_depth*3+93)-1:`VWidth*(`APPRam_depth*3+92)],data_in[`VWidth*(`APPRam_depth*2+93)-1:`VWidth*(`APPRam_depth*2+92)],data_in[`VWidth*(`APPRam_depth*1+93)-1:`VWidth*(`APPRam_depth*1+92)],data_in[`VWidth*(`APPRam_depth*0+93)-1:`VWidth*(`APPRam_depth*0+92)]};
			end
			93:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+94)-1:`VWidth*(`APPRam_depth*31+93)],data_in[`VWidth*(`APPRam_depth*30+94)-1:`VWidth*(`APPRam_depth*30+93)],data_in[`VWidth*(`APPRam_depth*29+94)-1:`VWidth*(`APPRam_depth*29+93)],data_in[`VWidth*(`APPRam_depth*28+94)-1:`VWidth*(`APPRam_depth*28+93)],data_in[`VWidth*(`APPRam_depth*27+94)-1:`VWidth*(`APPRam_depth*27+93)],data_in[`VWidth*(`APPRam_depth*26+94)-1:`VWidth*(`APPRam_depth*26+93)],data_in[`VWidth*(`APPRam_depth*25+94)-1:`VWidth*(`APPRam_depth*25+93)],data_in[`VWidth*(`APPRam_depth*24+94)-1:`VWidth*(`APPRam_depth*24+93)],data_in[`VWidth*(`APPRam_depth*23+94)-1:`VWidth*(`APPRam_depth*23+93)],data_in[`VWidth*(`APPRam_depth*22+94)-1:`VWidth*(`APPRam_depth*22+93)],data_in[`VWidth*(`APPRam_depth*21+94)-1:`VWidth*(`APPRam_depth*21+93)],data_in[`VWidth*(`APPRam_depth*20+94)-1:`VWidth*(`APPRam_depth*20+93)],data_in[`VWidth*(`APPRam_depth*19+94)-1:`VWidth*(`APPRam_depth*19+93)],data_in[`VWidth*(`APPRam_depth*18+94)-1:`VWidth*(`APPRam_depth*18+93)],data_in[`VWidth*(`APPRam_depth*17+94)-1:`VWidth*(`APPRam_depth*17+93)],data_in[`VWidth*(`APPRam_depth*16+94)-1:`VWidth*(`APPRam_depth*16+93)],data_in[`VWidth*(`APPRam_depth*15+94)-1:`VWidth*(`APPRam_depth*15+93)],data_in[`VWidth*(`APPRam_depth*14+94)-1:`VWidth*(`APPRam_depth*14+93)],data_in[`VWidth*(`APPRam_depth*13+94)-1:`VWidth*(`APPRam_depth*13+93)],data_in[`VWidth*(`APPRam_depth*12+94)-1:`VWidth*(`APPRam_depth*12+93)],data_in[`VWidth*(`APPRam_depth*11+94)-1:`VWidth*(`APPRam_depth*11+93)],data_in[`VWidth*(`APPRam_depth*10+94)-1:`VWidth*(`APPRam_depth*10+93)],data_in[`VWidth*(`APPRam_depth*9+94)-1:`VWidth*(`APPRam_depth*9+93)],data_in[`VWidth*(`APPRam_depth*8+94)-1:`VWidth*(`APPRam_depth*8+93)],data_in[`VWidth*(`APPRam_depth*7+94)-1:`VWidth*(`APPRam_depth*7+93)],data_in[`VWidth*(`APPRam_depth*6+94)-1:`VWidth*(`APPRam_depth*6+93)],data_in[`VWidth*(`APPRam_depth*5+94)-1:`VWidth*(`APPRam_depth*5+93)],data_in[`VWidth*(`APPRam_depth*4+94)-1:`VWidth*(`APPRam_depth*4+93)],data_in[`VWidth*(`APPRam_depth*3+94)-1:`VWidth*(`APPRam_depth*3+93)],data_in[`VWidth*(`APPRam_depth*2+94)-1:`VWidth*(`APPRam_depth*2+93)],data_in[`VWidth*(`APPRam_depth*1+94)-1:`VWidth*(`APPRam_depth*1+93)],data_in[`VWidth*(`APPRam_depth*0+94)-1:`VWidth*(`APPRam_depth*0+93)]};
			end
			94:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+95)-1:`VWidth*(`APPRam_depth*31+94)],data_in[`VWidth*(`APPRam_depth*30+95)-1:`VWidth*(`APPRam_depth*30+94)],data_in[`VWidth*(`APPRam_depth*29+95)-1:`VWidth*(`APPRam_depth*29+94)],data_in[`VWidth*(`APPRam_depth*28+95)-1:`VWidth*(`APPRam_depth*28+94)],data_in[`VWidth*(`APPRam_depth*27+95)-1:`VWidth*(`APPRam_depth*27+94)],data_in[`VWidth*(`APPRam_depth*26+95)-1:`VWidth*(`APPRam_depth*26+94)],data_in[`VWidth*(`APPRam_depth*25+95)-1:`VWidth*(`APPRam_depth*25+94)],data_in[`VWidth*(`APPRam_depth*24+95)-1:`VWidth*(`APPRam_depth*24+94)],data_in[`VWidth*(`APPRam_depth*23+95)-1:`VWidth*(`APPRam_depth*23+94)],data_in[`VWidth*(`APPRam_depth*22+95)-1:`VWidth*(`APPRam_depth*22+94)],data_in[`VWidth*(`APPRam_depth*21+95)-1:`VWidth*(`APPRam_depth*21+94)],data_in[`VWidth*(`APPRam_depth*20+95)-1:`VWidth*(`APPRam_depth*20+94)],data_in[`VWidth*(`APPRam_depth*19+95)-1:`VWidth*(`APPRam_depth*19+94)],data_in[`VWidth*(`APPRam_depth*18+95)-1:`VWidth*(`APPRam_depth*18+94)],data_in[`VWidth*(`APPRam_depth*17+95)-1:`VWidth*(`APPRam_depth*17+94)],data_in[`VWidth*(`APPRam_depth*16+95)-1:`VWidth*(`APPRam_depth*16+94)],data_in[`VWidth*(`APPRam_depth*15+95)-1:`VWidth*(`APPRam_depth*15+94)],data_in[`VWidth*(`APPRam_depth*14+95)-1:`VWidth*(`APPRam_depth*14+94)],data_in[`VWidth*(`APPRam_depth*13+95)-1:`VWidth*(`APPRam_depth*13+94)],data_in[`VWidth*(`APPRam_depth*12+95)-1:`VWidth*(`APPRam_depth*12+94)],data_in[`VWidth*(`APPRam_depth*11+95)-1:`VWidth*(`APPRam_depth*11+94)],data_in[`VWidth*(`APPRam_depth*10+95)-1:`VWidth*(`APPRam_depth*10+94)],data_in[`VWidth*(`APPRam_depth*9+95)-1:`VWidth*(`APPRam_depth*9+94)],data_in[`VWidth*(`APPRam_depth*8+95)-1:`VWidth*(`APPRam_depth*8+94)],data_in[`VWidth*(`APPRam_depth*7+95)-1:`VWidth*(`APPRam_depth*7+94)],data_in[`VWidth*(`APPRam_depth*6+95)-1:`VWidth*(`APPRam_depth*6+94)],data_in[`VWidth*(`APPRam_depth*5+95)-1:`VWidth*(`APPRam_depth*5+94)],data_in[`VWidth*(`APPRam_depth*4+95)-1:`VWidth*(`APPRam_depth*4+94)],data_in[`VWidth*(`APPRam_depth*3+95)-1:`VWidth*(`APPRam_depth*3+94)],data_in[`VWidth*(`APPRam_depth*2+95)-1:`VWidth*(`APPRam_depth*2+94)],data_in[`VWidth*(`APPRam_depth*1+95)-1:`VWidth*(`APPRam_depth*1+94)],data_in[`VWidth*(`APPRam_depth*0+95)-1:`VWidth*(`APPRam_depth*0+94)]};
			end
			95:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+96)-1:`VWidth*(`APPRam_depth*31+95)],data_in[`VWidth*(`APPRam_depth*30+96)-1:`VWidth*(`APPRam_depth*30+95)],data_in[`VWidth*(`APPRam_depth*29+96)-1:`VWidth*(`APPRam_depth*29+95)],data_in[`VWidth*(`APPRam_depth*28+96)-1:`VWidth*(`APPRam_depth*28+95)],data_in[`VWidth*(`APPRam_depth*27+96)-1:`VWidth*(`APPRam_depth*27+95)],data_in[`VWidth*(`APPRam_depth*26+96)-1:`VWidth*(`APPRam_depth*26+95)],data_in[`VWidth*(`APPRam_depth*25+96)-1:`VWidth*(`APPRam_depth*25+95)],data_in[`VWidth*(`APPRam_depth*24+96)-1:`VWidth*(`APPRam_depth*24+95)],data_in[`VWidth*(`APPRam_depth*23+96)-1:`VWidth*(`APPRam_depth*23+95)],data_in[`VWidth*(`APPRam_depth*22+96)-1:`VWidth*(`APPRam_depth*22+95)],data_in[`VWidth*(`APPRam_depth*21+96)-1:`VWidth*(`APPRam_depth*21+95)],data_in[`VWidth*(`APPRam_depth*20+96)-1:`VWidth*(`APPRam_depth*20+95)],data_in[`VWidth*(`APPRam_depth*19+96)-1:`VWidth*(`APPRam_depth*19+95)],data_in[`VWidth*(`APPRam_depth*18+96)-1:`VWidth*(`APPRam_depth*18+95)],data_in[`VWidth*(`APPRam_depth*17+96)-1:`VWidth*(`APPRam_depth*17+95)],data_in[`VWidth*(`APPRam_depth*16+96)-1:`VWidth*(`APPRam_depth*16+95)],data_in[`VWidth*(`APPRam_depth*15+96)-1:`VWidth*(`APPRam_depth*15+95)],data_in[`VWidth*(`APPRam_depth*14+96)-1:`VWidth*(`APPRam_depth*14+95)],data_in[`VWidth*(`APPRam_depth*13+96)-1:`VWidth*(`APPRam_depth*13+95)],data_in[`VWidth*(`APPRam_depth*12+96)-1:`VWidth*(`APPRam_depth*12+95)],data_in[`VWidth*(`APPRam_depth*11+96)-1:`VWidth*(`APPRam_depth*11+95)],data_in[`VWidth*(`APPRam_depth*10+96)-1:`VWidth*(`APPRam_depth*10+95)],data_in[`VWidth*(`APPRam_depth*9+96)-1:`VWidth*(`APPRam_depth*9+95)],data_in[`VWidth*(`APPRam_depth*8+96)-1:`VWidth*(`APPRam_depth*8+95)],data_in[`VWidth*(`APPRam_depth*7+96)-1:`VWidth*(`APPRam_depth*7+95)],data_in[`VWidth*(`APPRam_depth*6+96)-1:`VWidth*(`APPRam_depth*6+95)],data_in[`VWidth*(`APPRam_depth*5+96)-1:`VWidth*(`APPRam_depth*5+95)],data_in[`VWidth*(`APPRam_depth*4+96)-1:`VWidth*(`APPRam_depth*4+95)],data_in[`VWidth*(`APPRam_depth*3+96)-1:`VWidth*(`APPRam_depth*3+95)],data_in[`VWidth*(`APPRam_depth*2+96)-1:`VWidth*(`APPRam_depth*2+95)],data_in[`VWidth*(`APPRam_depth*1+96)-1:`VWidth*(`APPRam_depth*1+95)],data_in[`VWidth*(`APPRam_depth*0+96)-1:`VWidth*(`APPRam_depth*0+95)]};
			end
			96:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+97)-1:`VWidth*(`APPRam_depth*31+96)],data_in[`VWidth*(`APPRam_depth*30+97)-1:`VWidth*(`APPRam_depth*30+96)],data_in[`VWidth*(`APPRam_depth*29+97)-1:`VWidth*(`APPRam_depth*29+96)],data_in[`VWidth*(`APPRam_depth*28+97)-1:`VWidth*(`APPRam_depth*28+96)],data_in[`VWidth*(`APPRam_depth*27+97)-1:`VWidth*(`APPRam_depth*27+96)],data_in[`VWidth*(`APPRam_depth*26+97)-1:`VWidth*(`APPRam_depth*26+96)],data_in[`VWidth*(`APPRam_depth*25+97)-1:`VWidth*(`APPRam_depth*25+96)],data_in[`VWidth*(`APPRam_depth*24+97)-1:`VWidth*(`APPRam_depth*24+96)],data_in[`VWidth*(`APPRam_depth*23+97)-1:`VWidth*(`APPRam_depth*23+96)],data_in[`VWidth*(`APPRam_depth*22+97)-1:`VWidth*(`APPRam_depth*22+96)],data_in[`VWidth*(`APPRam_depth*21+97)-1:`VWidth*(`APPRam_depth*21+96)],data_in[`VWidth*(`APPRam_depth*20+97)-1:`VWidth*(`APPRam_depth*20+96)],data_in[`VWidth*(`APPRam_depth*19+97)-1:`VWidth*(`APPRam_depth*19+96)],data_in[`VWidth*(`APPRam_depth*18+97)-1:`VWidth*(`APPRam_depth*18+96)],data_in[`VWidth*(`APPRam_depth*17+97)-1:`VWidth*(`APPRam_depth*17+96)],data_in[`VWidth*(`APPRam_depth*16+97)-1:`VWidth*(`APPRam_depth*16+96)],data_in[`VWidth*(`APPRam_depth*15+97)-1:`VWidth*(`APPRam_depth*15+96)],data_in[`VWidth*(`APPRam_depth*14+97)-1:`VWidth*(`APPRam_depth*14+96)],data_in[`VWidth*(`APPRam_depth*13+97)-1:`VWidth*(`APPRam_depth*13+96)],data_in[`VWidth*(`APPRam_depth*12+97)-1:`VWidth*(`APPRam_depth*12+96)],data_in[`VWidth*(`APPRam_depth*11+97)-1:`VWidth*(`APPRam_depth*11+96)],data_in[`VWidth*(`APPRam_depth*10+97)-1:`VWidth*(`APPRam_depth*10+96)],data_in[`VWidth*(`APPRam_depth*9+97)-1:`VWidth*(`APPRam_depth*9+96)],data_in[`VWidth*(`APPRam_depth*8+97)-1:`VWidth*(`APPRam_depth*8+96)],data_in[`VWidth*(`APPRam_depth*7+97)-1:`VWidth*(`APPRam_depth*7+96)],data_in[`VWidth*(`APPRam_depth*6+97)-1:`VWidth*(`APPRam_depth*6+96)],data_in[`VWidth*(`APPRam_depth*5+97)-1:`VWidth*(`APPRam_depth*5+96)],data_in[`VWidth*(`APPRam_depth*4+97)-1:`VWidth*(`APPRam_depth*4+96)],data_in[`VWidth*(`APPRam_depth*3+97)-1:`VWidth*(`APPRam_depth*3+96)],data_in[`VWidth*(`APPRam_depth*2+97)-1:`VWidth*(`APPRam_depth*2+96)],data_in[`VWidth*(`APPRam_depth*1+97)-1:`VWidth*(`APPRam_depth*1+96)],data_in[`VWidth*(`APPRam_depth*0+97)-1:`VWidth*(`APPRam_depth*0+96)]};
			end
			97:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+98)-1:`VWidth*(`APPRam_depth*31+97)],data_in[`VWidth*(`APPRam_depth*30+98)-1:`VWidth*(`APPRam_depth*30+97)],data_in[`VWidth*(`APPRam_depth*29+98)-1:`VWidth*(`APPRam_depth*29+97)],data_in[`VWidth*(`APPRam_depth*28+98)-1:`VWidth*(`APPRam_depth*28+97)],data_in[`VWidth*(`APPRam_depth*27+98)-1:`VWidth*(`APPRam_depth*27+97)],data_in[`VWidth*(`APPRam_depth*26+98)-1:`VWidth*(`APPRam_depth*26+97)],data_in[`VWidth*(`APPRam_depth*25+98)-1:`VWidth*(`APPRam_depth*25+97)],data_in[`VWidth*(`APPRam_depth*24+98)-1:`VWidth*(`APPRam_depth*24+97)],data_in[`VWidth*(`APPRam_depth*23+98)-1:`VWidth*(`APPRam_depth*23+97)],data_in[`VWidth*(`APPRam_depth*22+98)-1:`VWidth*(`APPRam_depth*22+97)],data_in[`VWidth*(`APPRam_depth*21+98)-1:`VWidth*(`APPRam_depth*21+97)],data_in[`VWidth*(`APPRam_depth*20+98)-1:`VWidth*(`APPRam_depth*20+97)],data_in[`VWidth*(`APPRam_depth*19+98)-1:`VWidth*(`APPRam_depth*19+97)],data_in[`VWidth*(`APPRam_depth*18+98)-1:`VWidth*(`APPRam_depth*18+97)],data_in[`VWidth*(`APPRam_depth*17+98)-1:`VWidth*(`APPRam_depth*17+97)],data_in[`VWidth*(`APPRam_depth*16+98)-1:`VWidth*(`APPRam_depth*16+97)],data_in[`VWidth*(`APPRam_depth*15+98)-1:`VWidth*(`APPRam_depth*15+97)],data_in[`VWidth*(`APPRam_depth*14+98)-1:`VWidth*(`APPRam_depth*14+97)],data_in[`VWidth*(`APPRam_depth*13+98)-1:`VWidth*(`APPRam_depth*13+97)],data_in[`VWidth*(`APPRam_depth*12+98)-1:`VWidth*(`APPRam_depth*12+97)],data_in[`VWidth*(`APPRam_depth*11+98)-1:`VWidth*(`APPRam_depth*11+97)],data_in[`VWidth*(`APPRam_depth*10+98)-1:`VWidth*(`APPRam_depth*10+97)],data_in[`VWidth*(`APPRam_depth*9+98)-1:`VWidth*(`APPRam_depth*9+97)],data_in[`VWidth*(`APPRam_depth*8+98)-1:`VWidth*(`APPRam_depth*8+97)],data_in[`VWidth*(`APPRam_depth*7+98)-1:`VWidth*(`APPRam_depth*7+97)],data_in[`VWidth*(`APPRam_depth*6+98)-1:`VWidth*(`APPRam_depth*6+97)],data_in[`VWidth*(`APPRam_depth*5+98)-1:`VWidth*(`APPRam_depth*5+97)],data_in[`VWidth*(`APPRam_depth*4+98)-1:`VWidth*(`APPRam_depth*4+97)],data_in[`VWidth*(`APPRam_depth*3+98)-1:`VWidth*(`APPRam_depth*3+97)],data_in[`VWidth*(`APPRam_depth*2+98)-1:`VWidth*(`APPRam_depth*2+97)],data_in[`VWidth*(`APPRam_depth*1+98)-1:`VWidth*(`APPRam_depth*1+97)],data_in[`VWidth*(`APPRam_depth*0+98)-1:`VWidth*(`APPRam_depth*0+97)]};
			end
			98:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+99)-1:`VWidth*(`APPRam_depth*31+98)],data_in[`VWidth*(`APPRam_depth*30+99)-1:`VWidth*(`APPRam_depth*30+98)],data_in[`VWidth*(`APPRam_depth*29+99)-1:`VWidth*(`APPRam_depth*29+98)],data_in[`VWidth*(`APPRam_depth*28+99)-1:`VWidth*(`APPRam_depth*28+98)],data_in[`VWidth*(`APPRam_depth*27+99)-1:`VWidth*(`APPRam_depth*27+98)],data_in[`VWidth*(`APPRam_depth*26+99)-1:`VWidth*(`APPRam_depth*26+98)],data_in[`VWidth*(`APPRam_depth*25+99)-1:`VWidth*(`APPRam_depth*25+98)],data_in[`VWidth*(`APPRam_depth*24+99)-1:`VWidth*(`APPRam_depth*24+98)],data_in[`VWidth*(`APPRam_depth*23+99)-1:`VWidth*(`APPRam_depth*23+98)],data_in[`VWidth*(`APPRam_depth*22+99)-1:`VWidth*(`APPRam_depth*22+98)],data_in[`VWidth*(`APPRam_depth*21+99)-1:`VWidth*(`APPRam_depth*21+98)],data_in[`VWidth*(`APPRam_depth*20+99)-1:`VWidth*(`APPRam_depth*20+98)],data_in[`VWidth*(`APPRam_depth*19+99)-1:`VWidth*(`APPRam_depth*19+98)],data_in[`VWidth*(`APPRam_depth*18+99)-1:`VWidth*(`APPRam_depth*18+98)],data_in[`VWidth*(`APPRam_depth*17+99)-1:`VWidth*(`APPRam_depth*17+98)],data_in[`VWidth*(`APPRam_depth*16+99)-1:`VWidth*(`APPRam_depth*16+98)],data_in[`VWidth*(`APPRam_depth*15+99)-1:`VWidth*(`APPRam_depth*15+98)],data_in[`VWidth*(`APPRam_depth*14+99)-1:`VWidth*(`APPRam_depth*14+98)],data_in[`VWidth*(`APPRam_depth*13+99)-1:`VWidth*(`APPRam_depth*13+98)],data_in[`VWidth*(`APPRam_depth*12+99)-1:`VWidth*(`APPRam_depth*12+98)],data_in[`VWidth*(`APPRam_depth*11+99)-1:`VWidth*(`APPRam_depth*11+98)],data_in[`VWidth*(`APPRam_depth*10+99)-1:`VWidth*(`APPRam_depth*10+98)],data_in[`VWidth*(`APPRam_depth*9+99)-1:`VWidth*(`APPRam_depth*9+98)],data_in[`VWidth*(`APPRam_depth*8+99)-1:`VWidth*(`APPRam_depth*8+98)],data_in[`VWidth*(`APPRam_depth*7+99)-1:`VWidth*(`APPRam_depth*7+98)],data_in[`VWidth*(`APPRam_depth*6+99)-1:`VWidth*(`APPRam_depth*6+98)],data_in[`VWidth*(`APPRam_depth*5+99)-1:`VWidth*(`APPRam_depth*5+98)],data_in[`VWidth*(`APPRam_depth*4+99)-1:`VWidth*(`APPRam_depth*4+98)],data_in[`VWidth*(`APPRam_depth*3+99)-1:`VWidth*(`APPRam_depth*3+98)],data_in[`VWidth*(`APPRam_depth*2+99)-1:`VWidth*(`APPRam_depth*2+98)],data_in[`VWidth*(`APPRam_depth*1+99)-1:`VWidth*(`APPRam_depth*1+98)],data_in[`VWidth*(`APPRam_depth*0+99)-1:`VWidth*(`APPRam_depth*0+98)]};
			end
			99:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+100)-1:`VWidth*(`APPRam_depth*31+99)],data_in[`VWidth*(`APPRam_depth*30+100)-1:`VWidth*(`APPRam_depth*30+99)],data_in[`VWidth*(`APPRam_depth*29+100)-1:`VWidth*(`APPRam_depth*29+99)],data_in[`VWidth*(`APPRam_depth*28+100)-1:`VWidth*(`APPRam_depth*28+99)],data_in[`VWidth*(`APPRam_depth*27+100)-1:`VWidth*(`APPRam_depth*27+99)],data_in[`VWidth*(`APPRam_depth*26+100)-1:`VWidth*(`APPRam_depth*26+99)],data_in[`VWidth*(`APPRam_depth*25+100)-1:`VWidth*(`APPRam_depth*25+99)],data_in[`VWidth*(`APPRam_depth*24+100)-1:`VWidth*(`APPRam_depth*24+99)],data_in[`VWidth*(`APPRam_depth*23+100)-1:`VWidth*(`APPRam_depth*23+99)],data_in[`VWidth*(`APPRam_depth*22+100)-1:`VWidth*(`APPRam_depth*22+99)],data_in[`VWidth*(`APPRam_depth*21+100)-1:`VWidth*(`APPRam_depth*21+99)],data_in[`VWidth*(`APPRam_depth*20+100)-1:`VWidth*(`APPRam_depth*20+99)],data_in[`VWidth*(`APPRam_depth*19+100)-1:`VWidth*(`APPRam_depth*19+99)],data_in[`VWidth*(`APPRam_depth*18+100)-1:`VWidth*(`APPRam_depth*18+99)],data_in[`VWidth*(`APPRam_depth*17+100)-1:`VWidth*(`APPRam_depth*17+99)],data_in[`VWidth*(`APPRam_depth*16+100)-1:`VWidth*(`APPRam_depth*16+99)],data_in[`VWidth*(`APPRam_depth*15+100)-1:`VWidth*(`APPRam_depth*15+99)],data_in[`VWidth*(`APPRam_depth*14+100)-1:`VWidth*(`APPRam_depth*14+99)],data_in[`VWidth*(`APPRam_depth*13+100)-1:`VWidth*(`APPRam_depth*13+99)],data_in[`VWidth*(`APPRam_depth*12+100)-1:`VWidth*(`APPRam_depth*12+99)],data_in[`VWidth*(`APPRam_depth*11+100)-1:`VWidth*(`APPRam_depth*11+99)],data_in[`VWidth*(`APPRam_depth*10+100)-1:`VWidth*(`APPRam_depth*10+99)],data_in[`VWidth*(`APPRam_depth*9+100)-1:`VWidth*(`APPRam_depth*9+99)],data_in[`VWidth*(`APPRam_depth*8+100)-1:`VWidth*(`APPRam_depth*8+99)],data_in[`VWidth*(`APPRam_depth*7+100)-1:`VWidth*(`APPRam_depth*7+99)],data_in[`VWidth*(`APPRam_depth*6+100)-1:`VWidth*(`APPRam_depth*6+99)],data_in[`VWidth*(`APPRam_depth*5+100)-1:`VWidth*(`APPRam_depth*5+99)],data_in[`VWidth*(`APPRam_depth*4+100)-1:`VWidth*(`APPRam_depth*4+99)],data_in[`VWidth*(`APPRam_depth*3+100)-1:`VWidth*(`APPRam_depth*3+99)],data_in[`VWidth*(`APPRam_depth*2+100)-1:`VWidth*(`APPRam_depth*2+99)],data_in[`VWidth*(`APPRam_depth*1+100)-1:`VWidth*(`APPRam_depth*1+99)],data_in[`VWidth*(`APPRam_depth*0+100)-1:`VWidth*(`APPRam_depth*0+99)]};
			end
			100:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+101)-1:`VWidth*(`APPRam_depth*31+100)],data_in[`VWidth*(`APPRam_depth*30+101)-1:`VWidth*(`APPRam_depth*30+100)],data_in[`VWidth*(`APPRam_depth*29+101)-1:`VWidth*(`APPRam_depth*29+100)],data_in[`VWidth*(`APPRam_depth*28+101)-1:`VWidth*(`APPRam_depth*28+100)],data_in[`VWidth*(`APPRam_depth*27+101)-1:`VWidth*(`APPRam_depth*27+100)],data_in[`VWidth*(`APPRam_depth*26+101)-1:`VWidth*(`APPRam_depth*26+100)],data_in[`VWidth*(`APPRam_depth*25+101)-1:`VWidth*(`APPRam_depth*25+100)],data_in[`VWidth*(`APPRam_depth*24+101)-1:`VWidth*(`APPRam_depth*24+100)],data_in[`VWidth*(`APPRam_depth*23+101)-1:`VWidth*(`APPRam_depth*23+100)],data_in[`VWidth*(`APPRam_depth*22+101)-1:`VWidth*(`APPRam_depth*22+100)],data_in[`VWidth*(`APPRam_depth*21+101)-1:`VWidth*(`APPRam_depth*21+100)],data_in[`VWidth*(`APPRam_depth*20+101)-1:`VWidth*(`APPRam_depth*20+100)],data_in[`VWidth*(`APPRam_depth*19+101)-1:`VWidth*(`APPRam_depth*19+100)],data_in[`VWidth*(`APPRam_depth*18+101)-1:`VWidth*(`APPRam_depth*18+100)],data_in[`VWidth*(`APPRam_depth*17+101)-1:`VWidth*(`APPRam_depth*17+100)],data_in[`VWidth*(`APPRam_depth*16+101)-1:`VWidth*(`APPRam_depth*16+100)],data_in[`VWidth*(`APPRam_depth*15+101)-1:`VWidth*(`APPRam_depth*15+100)],data_in[`VWidth*(`APPRam_depth*14+101)-1:`VWidth*(`APPRam_depth*14+100)],data_in[`VWidth*(`APPRam_depth*13+101)-1:`VWidth*(`APPRam_depth*13+100)],data_in[`VWidth*(`APPRam_depth*12+101)-1:`VWidth*(`APPRam_depth*12+100)],data_in[`VWidth*(`APPRam_depth*11+101)-1:`VWidth*(`APPRam_depth*11+100)],data_in[`VWidth*(`APPRam_depth*10+101)-1:`VWidth*(`APPRam_depth*10+100)],data_in[`VWidth*(`APPRam_depth*9+101)-1:`VWidth*(`APPRam_depth*9+100)],data_in[`VWidth*(`APPRam_depth*8+101)-1:`VWidth*(`APPRam_depth*8+100)],data_in[`VWidth*(`APPRam_depth*7+101)-1:`VWidth*(`APPRam_depth*7+100)],data_in[`VWidth*(`APPRam_depth*6+101)-1:`VWidth*(`APPRam_depth*6+100)],data_in[`VWidth*(`APPRam_depth*5+101)-1:`VWidth*(`APPRam_depth*5+100)],data_in[`VWidth*(`APPRam_depth*4+101)-1:`VWidth*(`APPRam_depth*4+100)],data_in[`VWidth*(`APPRam_depth*3+101)-1:`VWidth*(`APPRam_depth*3+100)],data_in[`VWidth*(`APPRam_depth*2+101)-1:`VWidth*(`APPRam_depth*2+100)],data_in[`VWidth*(`APPRam_depth*1+101)-1:`VWidth*(`APPRam_depth*1+100)],data_in[`VWidth*(`APPRam_depth*0+101)-1:`VWidth*(`APPRam_depth*0+100)]};
			end
			101:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+102)-1:`VWidth*(`APPRam_depth*31+101)],data_in[`VWidth*(`APPRam_depth*30+102)-1:`VWidth*(`APPRam_depth*30+101)],data_in[`VWidth*(`APPRam_depth*29+102)-1:`VWidth*(`APPRam_depth*29+101)],data_in[`VWidth*(`APPRam_depth*28+102)-1:`VWidth*(`APPRam_depth*28+101)],data_in[`VWidth*(`APPRam_depth*27+102)-1:`VWidth*(`APPRam_depth*27+101)],data_in[`VWidth*(`APPRam_depth*26+102)-1:`VWidth*(`APPRam_depth*26+101)],data_in[`VWidth*(`APPRam_depth*25+102)-1:`VWidth*(`APPRam_depth*25+101)],data_in[`VWidth*(`APPRam_depth*24+102)-1:`VWidth*(`APPRam_depth*24+101)],data_in[`VWidth*(`APPRam_depth*23+102)-1:`VWidth*(`APPRam_depth*23+101)],data_in[`VWidth*(`APPRam_depth*22+102)-1:`VWidth*(`APPRam_depth*22+101)],data_in[`VWidth*(`APPRam_depth*21+102)-1:`VWidth*(`APPRam_depth*21+101)],data_in[`VWidth*(`APPRam_depth*20+102)-1:`VWidth*(`APPRam_depth*20+101)],data_in[`VWidth*(`APPRam_depth*19+102)-1:`VWidth*(`APPRam_depth*19+101)],data_in[`VWidth*(`APPRam_depth*18+102)-1:`VWidth*(`APPRam_depth*18+101)],data_in[`VWidth*(`APPRam_depth*17+102)-1:`VWidth*(`APPRam_depth*17+101)],data_in[`VWidth*(`APPRam_depth*16+102)-1:`VWidth*(`APPRam_depth*16+101)],data_in[`VWidth*(`APPRam_depth*15+102)-1:`VWidth*(`APPRam_depth*15+101)],data_in[`VWidth*(`APPRam_depth*14+102)-1:`VWidth*(`APPRam_depth*14+101)],data_in[`VWidth*(`APPRam_depth*13+102)-1:`VWidth*(`APPRam_depth*13+101)],data_in[`VWidth*(`APPRam_depth*12+102)-1:`VWidth*(`APPRam_depth*12+101)],data_in[`VWidth*(`APPRam_depth*11+102)-1:`VWidth*(`APPRam_depth*11+101)],data_in[`VWidth*(`APPRam_depth*10+102)-1:`VWidth*(`APPRam_depth*10+101)],data_in[`VWidth*(`APPRam_depth*9+102)-1:`VWidth*(`APPRam_depth*9+101)],data_in[`VWidth*(`APPRam_depth*8+102)-1:`VWidth*(`APPRam_depth*8+101)],data_in[`VWidth*(`APPRam_depth*7+102)-1:`VWidth*(`APPRam_depth*7+101)],data_in[`VWidth*(`APPRam_depth*6+102)-1:`VWidth*(`APPRam_depth*6+101)],data_in[`VWidth*(`APPRam_depth*5+102)-1:`VWidth*(`APPRam_depth*5+101)],data_in[`VWidth*(`APPRam_depth*4+102)-1:`VWidth*(`APPRam_depth*4+101)],data_in[`VWidth*(`APPRam_depth*3+102)-1:`VWidth*(`APPRam_depth*3+101)],data_in[`VWidth*(`APPRam_depth*2+102)-1:`VWidth*(`APPRam_depth*2+101)],data_in[`VWidth*(`APPRam_depth*1+102)-1:`VWidth*(`APPRam_depth*1+101)],data_in[`VWidth*(`APPRam_depth*0+102)-1:`VWidth*(`APPRam_depth*0+101)]};
			end
			102:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+103)-1:`VWidth*(`APPRam_depth*31+102)],data_in[`VWidth*(`APPRam_depth*30+103)-1:`VWidth*(`APPRam_depth*30+102)],data_in[`VWidth*(`APPRam_depth*29+103)-1:`VWidth*(`APPRam_depth*29+102)],data_in[`VWidth*(`APPRam_depth*28+103)-1:`VWidth*(`APPRam_depth*28+102)],data_in[`VWidth*(`APPRam_depth*27+103)-1:`VWidth*(`APPRam_depth*27+102)],data_in[`VWidth*(`APPRam_depth*26+103)-1:`VWidth*(`APPRam_depth*26+102)],data_in[`VWidth*(`APPRam_depth*25+103)-1:`VWidth*(`APPRam_depth*25+102)],data_in[`VWidth*(`APPRam_depth*24+103)-1:`VWidth*(`APPRam_depth*24+102)],data_in[`VWidth*(`APPRam_depth*23+103)-1:`VWidth*(`APPRam_depth*23+102)],data_in[`VWidth*(`APPRam_depth*22+103)-1:`VWidth*(`APPRam_depth*22+102)],data_in[`VWidth*(`APPRam_depth*21+103)-1:`VWidth*(`APPRam_depth*21+102)],data_in[`VWidth*(`APPRam_depth*20+103)-1:`VWidth*(`APPRam_depth*20+102)],data_in[`VWidth*(`APPRam_depth*19+103)-1:`VWidth*(`APPRam_depth*19+102)],data_in[`VWidth*(`APPRam_depth*18+103)-1:`VWidth*(`APPRam_depth*18+102)],data_in[`VWidth*(`APPRam_depth*17+103)-1:`VWidth*(`APPRam_depth*17+102)],data_in[`VWidth*(`APPRam_depth*16+103)-1:`VWidth*(`APPRam_depth*16+102)],data_in[`VWidth*(`APPRam_depth*15+103)-1:`VWidth*(`APPRam_depth*15+102)],data_in[`VWidth*(`APPRam_depth*14+103)-1:`VWidth*(`APPRam_depth*14+102)],data_in[`VWidth*(`APPRam_depth*13+103)-1:`VWidth*(`APPRam_depth*13+102)],data_in[`VWidth*(`APPRam_depth*12+103)-1:`VWidth*(`APPRam_depth*12+102)],data_in[`VWidth*(`APPRam_depth*11+103)-1:`VWidth*(`APPRam_depth*11+102)],data_in[`VWidth*(`APPRam_depth*10+103)-1:`VWidth*(`APPRam_depth*10+102)],data_in[`VWidth*(`APPRam_depth*9+103)-1:`VWidth*(`APPRam_depth*9+102)],data_in[`VWidth*(`APPRam_depth*8+103)-1:`VWidth*(`APPRam_depth*8+102)],data_in[`VWidth*(`APPRam_depth*7+103)-1:`VWidth*(`APPRam_depth*7+102)],data_in[`VWidth*(`APPRam_depth*6+103)-1:`VWidth*(`APPRam_depth*6+102)],data_in[`VWidth*(`APPRam_depth*5+103)-1:`VWidth*(`APPRam_depth*5+102)],data_in[`VWidth*(`APPRam_depth*4+103)-1:`VWidth*(`APPRam_depth*4+102)],data_in[`VWidth*(`APPRam_depth*3+103)-1:`VWidth*(`APPRam_depth*3+102)],data_in[`VWidth*(`APPRam_depth*2+103)-1:`VWidth*(`APPRam_depth*2+102)],data_in[`VWidth*(`APPRam_depth*1+103)-1:`VWidth*(`APPRam_depth*1+102)],data_in[`VWidth*(`APPRam_depth*0+103)-1:`VWidth*(`APPRam_depth*0+102)]};
			end
			103:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+104)-1:`VWidth*(`APPRam_depth*31+103)],data_in[`VWidth*(`APPRam_depth*30+104)-1:`VWidth*(`APPRam_depth*30+103)],data_in[`VWidth*(`APPRam_depth*29+104)-1:`VWidth*(`APPRam_depth*29+103)],data_in[`VWidth*(`APPRam_depth*28+104)-1:`VWidth*(`APPRam_depth*28+103)],data_in[`VWidth*(`APPRam_depth*27+104)-1:`VWidth*(`APPRam_depth*27+103)],data_in[`VWidth*(`APPRam_depth*26+104)-1:`VWidth*(`APPRam_depth*26+103)],data_in[`VWidth*(`APPRam_depth*25+104)-1:`VWidth*(`APPRam_depth*25+103)],data_in[`VWidth*(`APPRam_depth*24+104)-1:`VWidth*(`APPRam_depth*24+103)],data_in[`VWidth*(`APPRam_depth*23+104)-1:`VWidth*(`APPRam_depth*23+103)],data_in[`VWidth*(`APPRam_depth*22+104)-1:`VWidth*(`APPRam_depth*22+103)],data_in[`VWidth*(`APPRam_depth*21+104)-1:`VWidth*(`APPRam_depth*21+103)],data_in[`VWidth*(`APPRam_depth*20+104)-1:`VWidth*(`APPRam_depth*20+103)],data_in[`VWidth*(`APPRam_depth*19+104)-1:`VWidth*(`APPRam_depth*19+103)],data_in[`VWidth*(`APPRam_depth*18+104)-1:`VWidth*(`APPRam_depth*18+103)],data_in[`VWidth*(`APPRam_depth*17+104)-1:`VWidth*(`APPRam_depth*17+103)],data_in[`VWidth*(`APPRam_depth*16+104)-1:`VWidth*(`APPRam_depth*16+103)],data_in[`VWidth*(`APPRam_depth*15+104)-1:`VWidth*(`APPRam_depth*15+103)],data_in[`VWidth*(`APPRam_depth*14+104)-1:`VWidth*(`APPRam_depth*14+103)],data_in[`VWidth*(`APPRam_depth*13+104)-1:`VWidth*(`APPRam_depth*13+103)],data_in[`VWidth*(`APPRam_depth*12+104)-1:`VWidth*(`APPRam_depth*12+103)],data_in[`VWidth*(`APPRam_depth*11+104)-1:`VWidth*(`APPRam_depth*11+103)],data_in[`VWidth*(`APPRam_depth*10+104)-1:`VWidth*(`APPRam_depth*10+103)],data_in[`VWidth*(`APPRam_depth*9+104)-1:`VWidth*(`APPRam_depth*9+103)],data_in[`VWidth*(`APPRam_depth*8+104)-1:`VWidth*(`APPRam_depth*8+103)],data_in[`VWidth*(`APPRam_depth*7+104)-1:`VWidth*(`APPRam_depth*7+103)],data_in[`VWidth*(`APPRam_depth*6+104)-1:`VWidth*(`APPRam_depth*6+103)],data_in[`VWidth*(`APPRam_depth*5+104)-1:`VWidth*(`APPRam_depth*5+103)],data_in[`VWidth*(`APPRam_depth*4+104)-1:`VWidth*(`APPRam_depth*4+103)],data_in[`VWidth*(`APPRam_depth*3+104)-1:`VWidth*(`APPRam_depth*3+103)],data_in[`VWidth*(`APPRam_depth*2+104)-1:`VWidth*(`APPRam_depth*2+103)],data_in[`VWidth*(`APPRam_depth*1+104)-1:`VWidth*(`APPRam_depth*1+103)],data_in[`VWidth*(`APPRam_depth*0+104)-1:`VWidth*(`APPRam_depth*0+103)]};
			end
			104:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+105)-1:`VWidth*(`APPRam_depth*31+104)],data_in[`VWidth*(`APPRam_depth*30+105)-1:`VWidth*(`APPRam_depth*30+104)],data_in[`VWidth*(`APPRam_depth*29+105)-1:`VWidth*(`APPRam_depth*29+104)],data_in[`VWidth*(`APPRam_depth*28+105)-1:`VWidth*(`APPRam_depth*28+104)],data_in[`VWidth*(`APPRam_depth*27+105)-1:`VWidth*(`APPRam_depth*27+104)],data_in[`VWidth*(`APPRam_depth*26+105)-1:`VWidth*(`APPRam_depth*26+104)],data_in[`VWidth*(`APPRam_depth*25+105)-1:`VWidth*(`APPRam_depth*25+104)],data_in[`VWidth*(`APPRam_depth*24+105)-1:`VWidth*(`APPRam_depth*24+104)],data_in[`VWidth*(`APPRam_depth*23+105)-1:`VWidth*(`APPRam_depth*23+104)],data_in[`VWidth*(`APPRam_depth*22+105)-1:`VWidth*(`APPRam_depth*22+104)],data_in[`VWidth*(`APPRam_depth*21+105)-1:`VWidth*(`APPRam_depth*21+104)],data_in[`VWidth*(`APPRam_depth*20+105)-1:`VWidth*(`APPRam_depth*20+104)],data_in[`VWidth*(`APPRam_depth*19+105)-1:`VWidth*(`APPRam_depth*19+104)],data_in[`VWidth*(`APPRam_depth*18+105)-1:`VWidth*(`APPRam_depth*18+104)],data_in[`VWidth*(`APPRam_depth*17+105)-1:`VWidth*(`APPRam_depth*17+104)],data_in[`VWidth*(`APPRam_depth*16+105)-1:`VWidth*(`APPRam_depth*16+104)],data_in[`VWidth*(`APPRam_depth*15+105)-1:`VWidth*(`APPRam_depth*15+104)],data_in[`VWidth*(`APPRam_depth*14+105)-1:`VWidth*(`APPRam_depth*14+104)],data_in[`VWidth*(`APPRam_depth*13+105)-1:`VWidth*(`APPRam_depth*13+104)],data_in[`VWidth*(`APPRam_depth*12+105)-1:`VWidth*(`APPRam_depth*12+104)],data_in[`VWidth*(`APPRam_depth*11+105)-1:`VWidth*(`APPRam_depth*11+104)],data_in[`VWidth*(`APPRam_depth*10+105)-1:`VWidth*(`APPRam_depth*10+104)],data_in[`VWidth*(`APPRam_depth*9+105)-1:`VWidth*(`APPRam_depth*9+104)],data_in[`VWidth*(`APPRam_depth*8+105)-1:`VWidth*(`APPRam_depth*8+104)],data_in[`VWidth*(`APPRam_depth*7+105)-1:`VWidth*(`APPRam_depth*7+104)],data_in[`VWidth*(`APPRam_depth*6+105)-1:`VWidth*(`APPRam_depth*6+104)],data_in[`VWidth*(`APPRam_depth*5+105)-1:`VWidth*(`APPRam_depth*5+104)],data_in[`VWidth*(`APPRam_depth*4+105)-1:`VWidth*(`APPRam_depth*4+104)],data_in[`VWidth*(`APPRam_depth*3+105)-1:`VWidth*(`APPRam_depth*3+104)],data_in[`VWidth*(`APPRam_depth*2+105)-1:`VWidth*(`APPRam_depth*2+104)],data_in[`VWidth*(`APPRam_depth*1+105)-1:`VWidth*(`APPRam_depth*1+104)],data_in[`VWidth*(`APPRam_depth*0+105)-1:`VWidth*(`APPRam_depth*0+104)]};
			end
			105:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+106)-1:`VWidth*(`APPRam_depth*31+105)],data_in[`VWidth*(`APPRam_depth*30+106)-1:`VWidth*(`APPRam_depth*30+105)],data_in[`VWidth*(`APPRam_depth*29+106)-1:`VWidth*(`APPRam_depth*29+105)],data_in[`VWidth*(`APPRam_depth*28+106)-1:`VWidth*(`APPRam_depth*28+105)],data_in[`VWidth*(`APPRam_depth*27+106)-1:`VWidth*(`APPRam_depth*27+105)],data_in[`VWidth*(`APPRam_depth*26+106)-1:`VWidth*(`APPRam_depth*26+105)],data_in[`VWidth*(`APPRam_depth*25+106)-1:`VWidth*(`APPRam_depth*25+105)],data_in[`VWidth*(`APPRam_depth*24+106)-1:`VWidth*(`APPRam_depth*24+105)],data_in[`VWidth*(`APPRam_depth*23+106)-1:`VWidth*(`APPRam_depth*23+105)],data_in[`VWidth*(`APPRam_depth*22+106)-1:`VWidth*(`APPRam_depth*22+105)],data_in[`VWidth*(`APPRam_depth*21+106)-1:`VWidth*(`APPRam_depth*21+105)],data_in[`VWidth*(`APPRam_depth*20+106)-1:`VWidth*(`APPRam_depth*20+105)],data_in[`VWidth*(`APPRam_depth*19+106)-1:`VWidth*(`APPRam_depth*19+105)],data_in[`VWidth*(`APPRam_depth*18+106)-1:`VWidth*(`APPRam_depth*18+105)],data_in[`VWidth*(`APPRam_depth*17+106)-1:`VWidth*(`APPRam_depth*17+105)],data_in[`VWidth*(`APPRam_depth*16+106)-1:`VWidth*(`APPRam_depth*16+105)],data_in[`VWidth*(`APPRam_depth*15+106)-1:`VWidth*(`APPRam_depth*15+105)],data_in[`VWidth*(`APPRam_depth*14+106)-1:`VWidth*(`APPRam_depth*14+105)],data_in[`VWidth*(`APPRam_depth*13+106)-1:`VWidth*(`APPRam_depth*13+105)],data_in[`VWidth*(`APPRam_depth*12+106)-1:`VWidth*(`APPRam_depth*12+105)],data_in[`VWidth*(`APPRam_depth*11+106)-1:`VWidth*(`APPRam_depth*11+105)],data_in[`VWidth*(`APPRam_depth*10+106)-1:`VWidth*(`APPRam_depth*10+105)],data_in[`VWidth*(`APPRam_depth*9+106)-1:`VWidth*(`APPRam_depth*9+105)],data_in[`VWidth*(`APPRam_depth*8+106)-1:`VWidth*(`APPRam_depth*8+105)],data_in[`VWidth*(`APPRam_depth*7+106)-1:`VWidth*(`APPRam_depth*7+105)],data_in[`VWidth*(`APPRam_depth*6+106)-1:`VWidth*(`APPRam_depth*6+105)],data_in[`VWidth*(`APPRam_depth*5+106)-1:`VWidth*(`APPRam_depth*5+105)],data_in[`VWidth*(`APPRam_depth*4+106)-1:`VWidth*(`APPRam_depth*4+105)],data_in[`VWidth*(`APPRam_depth*3+106)-1:`VWidth*(`APPRam_depth*3+105)],data_in[`VWidth*(`APPRam_depth*2+106)-1:`VWidth*(`APPRam_depth*2+105)],data_in[`VWidth*(`APPRam_depth*1+106)-1:`VWidth*(`APPRam_depth*1+105)],data_in[`VWidth*(`APPRam_depth*0+106)-1:`VWidth*(`APPRam_depth*0+105)]};
			end
			106:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+107)-1:`VWidth*(`APPRam_depth*31+106)],data_in[`VWidth*(`APPRam_depth*30+107)-1:`VWidth*(`APPRam_depth*30+106)],data_in[`VWidth*(`APPRam_depth*29+107)-1:`VWidth*(`APPRam_depth*29+106)],data_in[`VWidth*(`APPRam_depth*28+107)-1:`VWidth*(`APPRam_depth*28+106)],data_in[`VWidth*(`APPRam_depth*27+107)-1:`VWidth*(`APPRam_depth*27+106)],data_in[`VWidth*(`APPRam_depth*26+107)-1:`VWidth*(`APPRam_depth*26+106)],data_in[`VWidth*(`APPRam_depth*25+107)-1:`VWidth*(`APPRam_depth*25+106)],data_in[`VWidth*(`APPRam_depth*24+107)-1:`VWidth*(`APPRam_depth*24+106)],data_in[`VWidth*(`APPRam_depth*23+107)-1:`VWidth*(`APPRam_depth*23+106)],data_in[`VWidth*(`APPRam_depth*22+107)-1:`VWidth*(`APPRam_depth*22+106)],data_in[`VWidth*(`APPRam_depth*21+107)-1:`VWidth*(`APPRam_depth*21+106)],data_in[`VWidth*(`APPRam_depth*20+107)-1:`VWidth*(`APPRam_depth*20+106)],data_in[`VWidth*(`APPRam_depth*19+107)-1:`VWidth*(`APPRam_depth*19+106)],data_in[`VWidth*(`APPRam_depth*18+107)-1:`VWidth*(`APPRam_depth*18+106)],data_in[`VWidth*(`APPRam_depth*17+107)-1:`VWidth*(`APPRam_depth*17+106)],data_in[`VWidth*(`APPRam_depth*16+107)-1:`VWidth*(`APPRam_depth*16+106)],data_in[`VWidth*(`APPRam_depth*15+107)-1:`VWidth*(`APPRam_depth*15+106)],data_in[`VWidth*(`APPRam_depth*14+107)-1:`VWidth*(`APPRam_depth*14+106)],data_in[`VWidth*(`APPRam_depth*13+107)-1:`VWidth*(`APPRam_depth*13+106)],data_in[`VWidth*(`APPRam_depth*12+107)-1:`VWidth*(`APPRam_depth*12+106)],data_in[`VWidth*(`APPRam_depth*11+107)-1:`VWidth*(`APPRam_depth*11+106)],data_in[`VWidth*(`APPRam_depth*10+107)-1:`VWidth*(`APPRam_depth*10+106)],data_in[`VWidth*(`APPRam_depth*9+107)-1:`VWidth*(`APPRam_depth*9+106)],data_in[`VWidth*(`APPRam_depth*8+107)-1:`VWidth*(`APPRam_depth*8+106)],data_in[`VWidth*(`APPRam_depth*7+107)-1:`VWidth*(`APPRam_depth*7+106)],data_in[`VWidth*(`APPRam_depth*6+107)-1:`VWidth*(`APPRam_depth*6+106)],data_in[`VWidth*(`APPRam_depth*5+107)-1:`VWidth*(`APPRam_depth*5+106)],data_in[`VWidth*(`APPRam_depth*4+107)-1:`VWidth*(`APPRam_depth*4+106)],data_in[`VWidth*(`APPRam_depth*3+107)-1:`VWidth*(`APPRam_depth*3+106)],data_in[`VWidth*(`APPRam_depth*2+107)-1:`VWidth*(`APPRam_depth*2+106)],data_in[`VWidth*(`APPRam_depth*1+107)-1:`VWidth*(`APPRam_depth*1+106)],data_in[`VWidth*(`APPRam_depth*0+107)-1:`VWidth*(`APPRam_depth*0+106)]};
			end
			107:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+108)-1:`VWidth*(`APPRam_depth*31+107)],data_in[`VWidth*(`APPRam_depth*30+108)-1:`VWidth*(`APPRam_depth*30+107)],data_in[`VWidth*(`APPRam_depth*29+108)-1:`VWidth*(`APPRam_depth*29+107)],data_in[`VWidth*(`APPRam_depth*28+108)-1:`VWidth*(`APPRam_depth*28+107)],data_in[`VWidth*(`APPRam_depth*27+108)-1:`VWidth*(`APPRam_depth*27+107)],data_in[`VWidth*(`APPRam_depth*26+108)-1:`VWidth*(`APPRam_depth*26+107)],data_in[`VWidth*(`APPRam_depth*25+108)-1:`VWidth*(`APPRam_depth*25+107)],data_in[`VWidth*(`APPRam_depth*24+108)-1:`VWidth*(`APPRam_depth*24+107)],data_in[`VWidth*(`APPRam_depth*23+108)-1:`VWidth*(`APPRam_depth*23+107)],data_in[`VWidth*(`APPRam_depth*22+108)-1:`VWidth*(`APPRam_depth*22+107)],data_in[`VWidth*(`APPRam_depth*21+108)-1:`VWidth*(`APPRam_depth*21+107)],data_in[`VWidth*(`APPRam_depth*20+108)-1:`VWidth*(`APPRam_depth*20+107)],data_in[`VWidth*(`APPRam_depth*19+108)-1:`VWidth*(`APPRam_depth*19+107)],data_in[`VWidth*(`APPRam_depth*18+108)-1:`VWidth*(`APPRam_depth*18+107)],data_in[`VWidth*(`APPRam_depth*17+108)-1:`VWidth*(`APPRam_depth*17+107)],data_in[`VWidth*(`APPRam_depth*16+108)-1:`VWidth*(`APPRam_depth*16+107)],data_in[`VWidth*(`APPRam_depth*15+108)-1:`VWidth*(`APPRam_depth*15+107)],data_in[`VWidth*(`APPRam_depth*14+108)-1:`VWidth*(`APPRam_depth*14+107)],data_in[`VWidth*(`APPRam_depth*13+108)-1:`VWidth*(`APPRam_depth*13+107)],data_in[`VWidth*(`APPRam_depth*12+108)-1:`VWidth*(`APPRam_depth*12+107)],data_in[`VWidth*(`APPRam_depth*11+108)-1:`VWidth*(`APPRam_depth*11+107)],data_in[`VWidth*(`APPRam_depth*10+108)-1:`VWidth*(`APPRam_depth*10+107)],data_in[`VWidth*(`APPRam_depth*9+108)-1:`VWidth*(`APPRam_depth*9+107)],data_in[`VWidth*(`APPRam_depth*8+108)-1:`VWidth*(`APPRam_depth*8+107)],data_in[`VWidth*(`APPRam_depth*7+108)-1:`VWidth*(`APPRam_depth*7+107)],data_in[`VWidth*(`APPRam_depth*6+108)-1:`VWidth*(`APPRam_depth*6+107)],data_in[`VWidth*(`APPRam_depth*5+108)-1:`VWidth*(`APPRam_depth*5+107)],data_in[`VWidth*(`APPRam_depth*4+108)-1:`VWidth*(`APPRam_depth*4+107)],data_in[`VWidth*(`APPRam_depth*3+108)-1:`VWidth*(`APPRam_depth*3+107)],data_in[`VWidth*(`APPRam_depth*2+108)-1:`VWidth*(`APPRam_depth*2+107)],data_in[`VWidth*(`APPRam_depth*1+108)-1:`VWidth*(`APPRam_depth*1+107)],data_in[`VWidth*(`APPRam_depth*0+108)-1:`VWidth*(`APPRam_depth*0+107)]};
			end
			108:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+109)-1:`VWidth*(`APPRam_depth*31+108)],data_in[`VWidth*(`APPRam_depth*30+109)-1:`VWidth*(`APPRam_depth*30+108)],data_in[`VWidth*(`APPRam_depth*29+109)-1:`VWidth*(`APPRam_depth*29+108)],data_in[`VWidth*(`APPRam_depth*28+109)-1:`VWidth*(`APPRam_depth*28+108)],data_in[`VWidth*(`APPRam_depth*27+109)-1:`VWidth*(`APPRam_depth*27+108)],data_in[`VWidth*(`APPRam_depth*26+109)-1:`VWidth*(`APPRam_depth*26+108)],data_in[`VWidth*(`APPRam_depth*25+109)-1:`VWidth*(`APPRam_depth*25+108)],data_in[`VWidth*(`APPRam_depth*24+109)-1:`VWidth*(`APPRam_depth*24+108)],data_in[`VWidth*(`APPRam_depth*23+109)-1:`VWidth*(`APPRam_depth*23+108)],data_in[`VWidth*(`APPRam_depth*22+109)-1:`VWidth*(`APPRam_depth*22+108)],data_in[`VWidth*(`APPRam_depth*21+109)-1:`VWidth*(`APPRam_depth*21+108)],data_in[`VWidth*(`APPRam_depth*20+109)-1:`VWidth*(`APPRam_depth*20+108)],data_in[`VWidth*(`APPRam_depth*19+109)-1:`VWidth*(`APPRam_depth*19+108)],data_in[`VWidth*(`APPRam_depth*18+109)-1:`VWidth*(`APPRam_depth*18+108)],data_in[`VWidth*(`APPRam_depth*17+109)-1:`VWidth*(`APPRam_depth*17+108)],data_in[`VWidth*(`APPRam_depth*16+109)-1:`VWidth*(`APPRam_depth*16+108)],data_in[`VWidth*(`APPRam_depth*15+109)-1:`VWidth*(`APPRam_depth*15+108)],data_in[`VWidth*(`APPRam_depth*14+109)-1:`VWidth*(`APPRam_depth*14+108)],data_in[`VWidth*(`APPRam_depth*13+109)-1:`VWidth*(`APPRam_depth*13+108)],data_in[`VWidth*(`APPRam_depth*12+109)-1:`VWidth*(`APPRam_depth*12+108)],data_in[`VWidth*(`APPRam_depth*11+109)-1:`VWidth*(`APPRam_depth*11+108)],data_in[`VWidth*(`APPRam_depth*10+109)-1:`VWidth*(`APPRam_depth*10+108)],data_in[`VWidth*(`APPRam_depth*9+109)-1:`VWidth*(`APPRam_depth*9+108)],data_in[`VWidth*(`APPRam_depth*8+109)-1:`VWidth*(`APPRam_depth*8+108)],data_in[`VWidth*(`APPRam_depth*7+109)-1:`VWidth*(`APPRam_depth*7+108)],data_in[`VWidth*(`APPRam_depth*6+109)-1:`VWidth*(`APPRam_depth*6+108)],data_in[`VWidth*(`APPRam_depth*5+109)-1:`VWidth*(`APPRam_depth*5+108)],data_in[`VWidth*(`APPRam_depth*4+109)-1:`VWidth*(`APPRam_depth*4+108)],data_in[`VWidth*(`APPRam_depth*3+109)-1:`VWidth*(`APPRam_depth*3+108)],data_in[`VWidth*(`APPRam_depth*2+109)-1:`VWidth*(`APPRam_depth*2+108)],data_in[`VWidth*(`APPRam_depth*1+109)-1:`VWidth*(`APPRam_depth*1+108)],data_in[`VWidth*(`APPRam_depth*0+109)-1:`VWidth*(`APPRam_depth*0+108)]};
			end
			109:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+110)-1:`VWidth*(`APPRam_depth*31+109)],data_in[`VWidth*(`APPRam_depth*30+110)-1:`VWidth*(`APPRam_depth*30+109)],data_in[`VWidth*(`APPRam_depth*29+110)-1:`VWidth*(`APPRam_depth*29+109)],data_in[`VWidth*(`APPRam_depth*28+110)-1:`VWidth*(`APPRam_depth*28+109)],data_in[`VWidth*(`APPRam_depth*27+110)-1:`VWidth*(`APPRam_depth*27+109)],data_in[`VWidth*(`APPRam_depth*26+110)-1:`VWidth*(`APPRam_depth*26+109)],data_in[`VWidth*(`APPRam_depth*25+110)-1:`VWidth*(`APPRam_depth*25+109)],data_in[`VWidth*(`APPRam_depth*24+110)-1:`VWidth*(`APPRam_depth*24+109)],data_in[`VWidth*(`APPRam_depth*23+110)-1:`VWidth*(`APPRam_depth*23+109)],data_in[`VWidth*(`APPRam_depth*22+110)-1:`VWidth*(`APPRam_depth*22+109)],data_in[`VWidth*(`APPRam_depth*21+110)-1:`VWidth*(`APPRam_depth*21+109)],data_in[`VWidth*(`APPRam_depth*20+110)-1:`VWidth*(`APPRam_depth*20+109)],data_in[`VWidth*(`APPRam_depth*19+110)-1:`VWidth*(`APPRam_depth*19+109)],data_in[`VWidth*(`APPRam_depth*18+110)-1:`VWidth*(`APPRam_depth*18+109)],data_in[`VWidth*(`APPRam_depth*17+110)-1:`VWidth*(`APPRam_depth*17+109)],data_in[`VWidth*(`APPRam_depth*16+110)-1:`VWidth*(`APPRam_depth*16+109)],data_in[`VWidth*(`APPRam_depth*15+110)-1:`VWidth*(`APPRam_depth*15+109)],data_in[`VWidth*(`APPRam_depth*14+110)-1:`VWidth*(`APPRam_depth*14+109)],data_in[`VWidth*(`APPRam_depth*13+110)-1:`VWidth*(`APPRam_depth*13+109)],data_in[`VWidth*(`APPRam_depth*12+110)-1:`VWidth*(`APPRam_depth*12+109)],data_in[`VWidth*(`APPRam_depth*11+110)-1:`VWidth*(`APPRam_depth*11+109)],data_in[`VWidth*(`APPRam_depth*10+110)-1:`VWidth*(`APPRam_depth*10+109)],data_in[`VWidth*(`APPRam_depth*9+110)-1:`VWidth*(`APPRam_depth*9+109)],data_in[`VWidth*(`APPRam_depth*8+110)-1:`VWidth*(`APPRam_depth*8+109)],data_in[`VWidth*(`APPRam_depth*7+110)-1:`VWidth*(`APPRam_depth*7+109)],data_in[`VWidth*(`APPRam_depth*6+110)-1:`VWidth*(`APPRam_depth*6+109)],data_in[`VWidth*(`APPRam_depth*5+110)-1:`VWidth*(`APPRam_depth*5+109)],data_in[`VWidth*(`APPRam_depth*4+110)-1:`VWidth*(`APPRam_depth*4+109)],data_in[`VWidth*(`APPRam_depth*3+110)-1:`VWidth*(`APPRam_depth*3+109)],data_in[`VWidth*(`APPRam_depth*2+110)-1:`VWidth*(`APPRam_depth*2+109)],data_in[`VWidth*(`APPRam_depth*1+110)-1:`VWidth*(`APPRam_depth*1+109)],data_in[`VWidth*(`APPRam_depth*0+110)-1:`VWidth*(`APPRam_depth*0+109)]};
			end
			110:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+111)-1:`VWidth*(`APPRam_depth*31+110)],data_in[`VWidth*(`APPRam_depth*30+111)-1:`VWidth*(`APPRam_depth*30+110)],data_in[`VWidth*(`APPRam_depth*29+111)-1:`VWidth*(`APPRam_depth*29+110)],data_in[`VWidth*(`APPRam_depth*28+111)-1:`VWidth*(`APPRam_depth*28+110)],data_in[`VWidth*(`APPRam_depth*27+111)-1:`VWidth*(`APPRam_depth*27+110)],data_in[`VWidth*(`APPRam_depth*26+111)-1:`VWidth*(`APPRam_depth*26+110)],data_in[`VWidth*(`APPRam_depth*25+111)-1:`VWidth*(`APPRam_depth*25+110)],data_in[`VWidth*(`APPRam_depth*24+111)-1:`VWidth*(`APPRam_depth*24+110)],data_in[`VWidth*(`APPRam_depth*23+111)-1:`VWidth*(`APPRam_depth*23+110)],data_in[`VWidth*(`APPRam_depth*22+111)-1:`VWidth*(`APPRam_depth*22+110)],data_in[`VWidth*(`APPRam_depth*21+111)-1:`VWidth*(`APPRam_depth*21+110)],data_in[`VWidth*(`APPRam_depth*20+111)-1:`VWidth*(`APPRam_depth*20+110)],data_in[`VWidth*(`APPRam_depth*19+111)-1:`VWidth*(`APPRam_depth*19+110)],data_in[`VWidth*(`APPRam_depth*18+111)-1:`VWidth*(`APPRam_depth*18+110)],data_in[`VWidth*(`APPRam_depth*17+111)-1:`VWidth*(`APPRam_depth*17+110)],data_in[`VWidth*(`APPRam_depth*16+111)-1:`VWidth*(`APPRam_depth*16+110)],data_in[`VWidth*(`APPRam_depth*15+111)-1:`VWidth*(`APPRam_depth*15+110)],data_in[`VWidth*(`APPRam_depth*14+111)-1:`VWidth*(`APPRam_depth*14+110)],data_in[`VWidth*(`APPRam_depth*13+111)-1:`VWidth*(`APPRam_depth*13+110)],data_in[`VWidth*(`APPRam_depth*12+111)-1:`VWidth*(`APPRam_depth*12+110)],data_in[`VWidth*(`APPRam_depth*11+111)-1:`VWidth*(`APPRam_depth*11+110)],data_in[`VWidth*(`APPRam_depth*10+111)-1:`VWidth*(`APPRam_depth*10+110)],data_in[`VWidth*(`APPRam_depth*9+111)-1:`VWidth*(`APPRam_depth*9+110)],data_in[`VWidth*(`APPRam_depth*8+111)-1:`VWidth*(`APPRam_depth*8+110)],data_in[`VWidth*(`APPRam_depth*7+111)-1:`VWidth*(`APPRam_depth*7+110)],data_in[`VWidth*(`APPRam_depth*6+111)-1:`VWidth*(`APPRam_depth*6+110)],data_in[`VWidth*(`APPRam_depth*5+111)-1:`VWidth*(`APPRam_depth*5+110)],data_in[`VWidth*(`APPRam_depth*4+111)-1:`VWidth*(`APPRam_depth*4+110)],data_in[`VWidth*(`APPRam_depth*3+111)-1:`VWidth*(`APPRam_depth*3+110)],data_in[`VWidth*(`APPRam_depth*2+111)-1:`VWidth*(`APPRam_depth*2+110)],data_in[`VWidth*(`APPRam_depth*1+111)-1:`VWidth*(`APPRam_depth*1+110)],data_in[`VWidth*(`APPRam_depth*0+111)-1:`VWidth*(`APPRam_depth*0+110)]};
			end
			111:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+112)-1:`VWidth*(`APPRam_depth*31+111)],data_in[`VWidth*(`APPRam_depth*30+112)-1:`VWidth*(`APPRam_depth*30+111)],data_in[`VWidth*(`APPRam_depth*29+112)-1:`VWidth*(`APPRam_depth*29+111)],data_in[`VWidth*(`APPRam_depth*28+112)-1:`VWidth*(`APPRam_depth*28+111)],data_in[`VWidth*(`APPRam_depth*27+112)-1:`VWidth*(`APPRam_depth*27+111)],data_in[`VWidth*(`APPRam_depth*26+112)-1:`VWidth*(`APPRam_depth*26+111)],data_in[`VWidth*(`APPRam_depth*25+112)-1:`VWidth*(`APPRam_depth*25+111)],data_in[`VWidth*(`APPRam_depth*24+112)-1:`VWidth*(`APPRam_depth*24+111)],data_in[`VWidth*(`APPRam_depth*23+112)-1:`VWidth*(`APPRam_depth*23+111)],data_in[`VWidth*(`APPRam_depth*22+112)-1:`VWidth*(`APPRam_depth*22+111)],data_in[`VWidth*(`APPRam_depth*21+112)-1:`VWidth*(`APPRam_depth*21+111)],data_in[`VWidth*(`APPRam_depth*20+112)-1:`VWidth*(`APPRam_depth*20+111)],data_in[`VWidth*(`APPRam_depth*19+112)-1:`VWidth*(`APPRam_depth*19+111)],data_in[`VWidth*(`APPRam_depth*18+112)-1:`VWidth*(`APPRam_depth*18+111)],data_in[`VWidth*(`APPRam_depth*17+112)-1:`VWidth*(`APPRam_depth*17+111)],data_in[`VWidth*(`APPRam_depth*16+112)-1:`VWidth*(`APPRam_depth*16+111)],data_in[`VWidth*(`APPRam_depth*15+112)-1:`VWidth*(`APPRam_depth*15+111)],data_in[`VWidth*(`APPRam_depth*14+112)-1:`VWidth*(`APPRam_depth*14+111)],data_in[`VWidth*(`APPRam_depth*13+112)-1:`VWidth*(`APPRam_depth*13+111)],data_in[`VWidth*(`APPRam_depth*12+112)-1:`VWidth*(`APPRam_depth*12+111)],data_in[`VWidth*(`APPRam_depth*11+112)-1:`VWidth*(`APPRam_depth*11+111)],data_in[`VWidth*(`APPRam_depth*10+112)-1:`VWidth*(`APPRam_depth*10+111)],data_in[`VWidth*(`APPRam_depth*9+112)-1:`VWidth*(`APPRam_depth*9+111)],data_in[`VWidth*(`APPRam_depth*8+112)-1:`VWidth*(`APPRam_depth*8+111)],data_in[`VWidth*(`APPRam_depth*7+112)-1:`VWidth*(`APPRam_depth*7+111)],data_in[`VWidth*(`APPRam_depth*6+112)-1:`VWidth*(`APPRam_depth*6+111)],data_in[`VWidth*(`APPRam_depth*5+112)-1:`VWidth*(`APPRam_depth*5+111)],data_in[`VWidth*(`APPRam_depth*4+112)-1:`VWidth*(`APPRam_depth*4+111)],data_in[`VWidth*(`APPRam_depth*3+112)-1:`VWidth*(`APPRam_depth*3+111)],data_in[`VWidth*(`APPRam_depth*2+112)-1:`VWidth*(`APPRam_depth*2+111)],data_in[`VWidth*(`APPRam_depth*1+112)-1:`VWidth*(`APPRam_depth*1+111)],data_in[`VWidth*(`APPRam_depth*0+112)-1:`VWidth*(`APPRam_depth*0+111)]};
			end
			112:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+113)-1:`VWidth*(`APPRam_depth*31+112)],data_in[`VWidth*(`APPRam_depth*30+113)-1:`VWidth*(`APPRam_depth*30+112)],data_in[`VWidth*(`APPRam_depth*29+113)-1:`VWidth*(`APPRam_depth*29+112)],data_in[`VWidth*(`APPRam_depth*28+113)-1:`VWidth*(`APPRam_depth*28+112)],data_in[`VWidth*(`APPRam_depth*27+113)-1:`VWidth*(`APPRam_depth*27+112)],data_in[`VWidth*(`APPRam_depth*26+113)-1:`VWidth*(`APPRam_depth*26+112)],data_in[`VWidth*(`APPRam_depth*25+113)-1:`VWidth*(`APPRam_depth*25+112)],data_in[`VWidth*(`APPRam_depth*24+113)-1:`VWidth*(`APPRam_depth*24+112)],data_in[`VWidth*(`APPRam_depth*23+113)-1:`VWidth*(`APPRam_depth*23+112)],data_in[`VWidth*(`APPRam_depth*22+113)-1:`VWidth*(`APPRam_depth*22+112)],data_in[`VWidth*(`APPRam_depth*21+113)-1:`VWidth*(`APPRam_depth*21+112)],data_in[`VWidth*(`APPRam_depth*20+113)-1:`VWidth*(`APPRam_depth*20+112)],data_in[`VWidth*(`APPRam_depth*19+113)-1:`VWidth*(`APPRam_depth*19+112)],data_in[`VWidth*(`APPRam_depth*18+113)-1:`VWidth*(`APPRam_depth*18+112)],data_in[`VWidth*(`APPRam_depth*17+113)-1:`VWidth*(`APPRam_depth*17+112)],data_in[`VWidth*(`APPRam_depth*16+113)-1:`VWidth*(`APPRam_depth*16+112)],data_in[`VWidth*(`APPRam_depth*15+113)-1:`VWidth*(`APPRam_depth*15+112)],data_in[`VWidth*(`APPRam_depth*14+113)-1:`VWidth*(`APPRam_depth*14+112)],data_in[`VWidth*(`APPRam_depth*13+113)-1:`VWidth*(`APPRam_depth*13+112)],data_in[`VWidth*(`APPRam_depth*12+113)-1:`VWidth*(`APPRam_depth*12+112)],data_in[`VWidth*(`APPRam_depth*11+113)-1:`VWidth*(`APPRam_depth*11+112)],data_in[`VWidth*(`APPRam_depth*10+113)-1:`VWidth*(`APPRam_depth*10+112)],data_in[`VWidth*(`APPRam_depth*9+113)-1:`VWidth*(`APPRam_depth*9+112)],data_in[`VWidth*(`APPRam_depth*8+113)-1:`VWidth*(`APPRam_depth*8+112)],data_in[`VWidth*(`APPRam_depth*7+113)-1:`VWidth*(`APPRam_depth*7+112)],data_in[`VWidth*(`APPRam_depth*6+113)-1:`VWidth*(`APPRam_depth*6+112)],data_in[`VWidth*(`APPRam_depth*5+113)-1:`VWidth*(`APPRam_depth*5+112)],data_in[`VWidth*(`APPRam_depth*4+113)-1:`VWidth*(`APPRam_depth*4+112)],data_in[`VWidth*(`APPRam_depth*3+113)-1:`VWidth*(`APPRam_depth*3+112)],data_in[`VWidth*(`APPRam_depth*2+113)-1:`VWidth*(`APPRam_depth*2+112)],data_in[`VWidth*(`APPRam_depth*1+113)-1:`VWidth*(`APPRam_depth*1+112)],data_in[`VWidth*(`APPRam_depth*0+113)-1:`VWidth*(`APPRam_depth*0+112)]};
			end
			113:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+114)-1:`VWidth*(`APPRam_depth*31+113)],data_in[`VWidth*(`APPRam_depth*30+114)-1:`VWidth*(`APPRam_depth*30+113)],data_in[`VWidth*(`APPRam_depth*29+114)-1:`VWidth*(`APPRam_depth*29+113)],data_in[`VWidth*(`APPRam_depth*28+114)-1:`VWidth*(`APPRam_depth*28+113)],data_in[`VWidth*(`APPRam_depth*27+114)-1:`VWidth*(`APPRam_depth*27+113)],data_in[`VWidth*(`APPRam_depth*26+114)-1:`VWidth*(`APPRam_depth*26+113)],data_in[`VWidth*(`APPRam_depth*25+114)-1:`VWidth*(`APPRam_depth*25+113)],data_in[`VWidth*(`APPRam_depth*24+114)-1:`VWidth*(`APPRam_depth*24+113)],data_in[`VWidth*(`APPRam_depth*23+114)-1:`VWidth*(`APPRam_depth*23+113)],data_in[`VWidth*(`APPRam_depth*22+114)-1:`VWidth*(`APPRam_depth*22+113)],data_in[`VWidth*(`APPRam_depth*21+114)-1:`VWidth*(`APPRam_depth*21+113)],data_in[`VWidth*(`APPRam_depth*20+114)-1:`VWidth*(`APPRam_depth*20+113)],data_in[`VWidth*(`APPRam_depth*19+114)-1:`VWidth*(`APPRam_depth*19+113)],data_in[`VWidth*(`APPRam_depth*18+114)-1:`VWidth*(`APPRam_depth*18+113)],data_in[`VWidth*(`APPRam_depth*17+114)-1:`VWidth*(`APPRam_depth*17+113)],data_in[`VWidth*(`APPRam_depth*16+114)-1:`VWidth*(`APPRam_depth*16+113)],data_in[`VWidth*(`APPRam_depth*15+114)-1:`VWidth*(`APPRam_depth*15+113)],data_in[`VWidth*(`APPRam_depth*14+114)-1:`VWidth*(`APPRam_depth*14+113)],data_in[`VWidth*(`APPRam_depth*13+114)-1:`VWidth*(`APPRam_depth*13+113)],data_in[`VWidth*(`APPRam_depth*12+114)-1:`VWidth*(`APPRam_depth*12+113)],data_in[`VWidth*(`APPRam_depth*11+114)-1:`VWidth*(`APPRam_depth*11+113)],data_in[`VWidth*(`APPRam_depth*10+114)-1:`VWidth*(`APPRam_depth*10+113)],data_in[`VWidth*(`APPRam_depth*9+114)-1:`VWidth*(`APPRam_depth*9+113)],data_in[`VWidth*(`APPRam_depth*8+114)-1:`VWidth*(`APPRam_depth*8+113)],data_in[`VWidth*(`APPRam_depth*7+114)-1:`VWidth*(`APPRam_depth*7+113)],data_in[`VWidth*(`APPRam_depth*6+114)-1:`VWidth*(`APPRam_depth*6+113)],data_in[`VWidth*(`APPRam_depth*5+114)-1:`VWidth*(`APPRam_depth*5+113)],data_in[`VWidth*(`APPRam_depth*4+114)-1:`VWidth*(`APPRam_depth*4+113)],data_in[`VWidth*(`APPRam_depth*3+114)-1:`VWidth*(`APPRam_depth*3+113)],data_in[`VWidth*(`APPRam_depth*2+114)-1:`VWidth*(`APPRam_depth*2+113)],data_in[`VWidth*(`APPRam_depth*1+114)-1:`VWidth*(`APPRam_depth*1+113)],data_in[`VWidth*(`APPRam_depth*0+114)-1:`VWidth*(`APPRam_depth*0+113)]};
			end
			114:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+115)-1:`VWidth*(`APPRam_depth*31+114)],data_in[`VWidth*(`APPRam_depth*30+115)-1:`VWidth*(`APPRam_depth*30+114)],data_in[`VWidth*(`APPRam_depth*29+115)-1:`VWidth*(`APPRam_depth*29+114)],data_in[`VWidth*(`APPRam_depth*28+115)-1:`VWidth*(`APPRam_depth*28+114)],data_in[`VWidth*(`APPRam_depth*27+115)-1:`VWidth*(`APPRam_depth*27+114)],data_in[`VWidth*(`APPRam_depth*26+115)-1:`VWidth*(`APPRam_depth*26+114)],data_in[`VWidth*(`APPRam_depth*25+115)-1:`VWidth*(`APPRam_depth*25+114)],data_in[`VWidth*(`APPRam_depth*24+115)-1:`VWidth*(`APPRam_depth*24+114)],data_in[`VWidth*(`APPRam_depth*23+115)-1:`VWidth*(`APPRam_depth*23+114)],data_in[`VWidth*(`APPRam_depth*22+115)-1:`VWidth*(`APPRam_depth*22+114)],data_in[`VWidth*(`APPRam_depth*21+115)-1:`VWidth*(`APPRam_depth*21+114)],data_in[`VWidth*(`APPRam_depth*20+115)-1:`VWidth*(`APPRam_depth*20+114)],data_in[`VWidth*(`APPRam_depth*19+115)-1:`VWidth*(`APPRam_depth*19+114)],data_in[`VWidth*(`APPRam_depth*18+115)-1:`VWidth*(`APPRam_depth*18+114)],data_in[`VWidth*(`APPRam_depth*17+115)-1:`VWidth*(`APPRam_depth*17+114)],data_in[`VWidth*(`APPRam_depth*16+115)-1:`VWidth*(`APPRam_depth*16+114)],data_in[`VWidth*(`APPRam_depth*15+115)-1:`VWidth*(`APPRam_depth*15+114)],data_in[`VWidth*(`APPRam_depth*14+115)-1:`VWidth*(`APPRam_depth*14+114)],data_in[`VWidth*(`APPRam_depth*13+115)-1:`VWidth*(`APPRam_depth*13+114)],data_in[`VWidth*(`APPRam_depth*12+115)-1:`VWidth*(`APPRam_depth*12+114)],data_in[`VWidth*(`APPRam_depth*11+115)-1:`VWidth*(`APPRam_depth*11+114)],data_in[`VWidth*(`APPRam_depth*10+115)-1:`VWidth*(`APPRam_depth*10+114)],data_in[`VWidth*(`APPRam_depth*9+115)-1:`VWidth*(`APPRam_depth*9+114)],data_in[`VWidth*(`APPRam_depth*8+115)-1:`VWidth*(`APPRam_depth*8+114)],data_in[`VWidth*(`APPRam_depth*7+115)-1:`VWidth*(`APPRam_depth*7+114)],data_in[`VWidth*(`APPRam_depth*6+115)-1:`VWidth*(`APPRam_depth*6+114)],data_in[`VWidth*(`APPRam_depth*5+115)-1:`VWidth*(`APPRam_depth*5+114)],data_in[`VWidth*(`APPRam_depth*4+115)-1:`VWidth*(`APPRam_depth*4+114)],data_in[`VWidth*(`APPRam_depth*3+115)-1:`VWidth*(`APPRam_depth*3+114)],data_in[`VWidth*(`APPRam_depth*2+115)-1:`VWidth*(`APPRam_depth*2+114)],data_in[`VWidth*(`APPRam_depth*1+115)-1:`VWidth*(`APPRam_depth*1+114)],data_in[`VWidth*(`APPRam_depth*0+115)-1:`VWidth*(`APPRam_depth*0+114)]};
			end
			115:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+116)-1:`VWidth*(`APPRam_depth*31+115)],data_in[`VWidth*(`APPRam_depth*30+116)-1:`VWidth*(`APPRam_depth*30+115)],data_in[`VWidth*(`APPRam_depth*29+116)-1:`VWidth*(`APPRam_depth*29+115)],data_in[`VWidth*(`APPRam_depth*28+116)-1:`VWidth*(`APPRam_depth*28+115)],data_in[`VWidth*(`APPRam_depth*27+116)-1:`VWidth*(`APPRam_depth*27+115)],data_in[`VWidth*(`APPRam_depth*26+116)-1:`VWidth*(`APPRam_depth*26+115)],data_in[`VWidth*(`APPRam_depth*25+116)-1:`VWidth*(`APPRam_depth*25+115)],data_in[`VWidth*(`APPRam_depth*24+116)-1:`VWidth*(`APPRam_depth*24+115)],data_in[`VWidth*(`APPRam_depth*23+116)-1:`VWidth*(`APPRam_depth*23+115)],data_in[`VWidth*(`APPRam_depth*22+116)-1:`VWidth*(`APPRam_depth*22+115)],data_in[`VWidth*(`APPRam_depth*21+116)-1:`VWidth*(`APPRam_depth*21+115)],data_in[`VWidth*(`APPRam_depth*20+116)-1:`VWidth*(`APPRam_depth*20+115)],data_in[`VWidth*(`APPRam_depth*19+116)-1:`VWidth*(`APPRam_depth*19+115)],data_in[`VWidth*(`APPRam_depth*18+116)-1:`VWidth*(`APPRam_depth*18+115)],data_in[`VWidth*(`APPRam_depth*17+116)-1:`VWidth*(`APPRam_depth*17+115)],data_in[`VWidth*(`APPRam_depth*16+116)-1:`VWidth*(`APPRam_depth*16+115)],data_in[`VWidth*(`APPRam_depth*15+116)-1:`VWidth*(`APPRam_depth*15+115)],data_in[`VWidth*(`APPRam_depth*14+116)-1:`VWidth*(`APPRam_depth*14+115)],data_in[`VWidth*(`APPRam_depth*13+116)-1:`VWidth*(`APPRam_depth*13+115)],data_in[`VWidth*(`APPRam_depth*12+116)-1:`VWidth*(`APPRam_depth*12+115)],data_in[`VWidth*(`APPRam_depth*11+116)-1:`VWidth*(`APPRam_depth*11+115)],data_in[`VWidth*(`APPRam_depth*10+116)-1:`VWidth*(`APPRam_depth*10+115)],data_in[`VWidth*(`APPRam_depth*9+116)-1:`VWidth*(`APPRam_depth*9+115)],data_in[`VWidth*(`APPRam_depth*8+116)-1:`VWidth*(`APPRam_depth*8+115)],data_in[`VWidth*(`APPRam_depth*7+116)-1:`VWidth*(`APPRam_depth*7+115)],data_in[`VWidth*(`APPRam_depth*6+116)-1:`VWidth*(`APPRam_depth*6+115)],data_in[`VWidth*(`APPRam_depth*5+116)-1:`VWidth*(`APPRam_depth*5+115)],data_in[`VWidth*(`APPRam_depth*4+116)-1:`VWidth*(`APPRam_depth*4+115)],data_in[`VWidth*(`APPRam_depth*3+116)-1:`VWidth*(`APPRam_depth*3+115)],data_in[`VWidth*(`APPRam_depth*2+116)-1:`VWidth*(`APPRam_depth*2+115)],data_in[`VWidth*(`APPRam_depth*1+116)-1:`VWidth*(`APPRam_depth*1+115)],data_in[`VWidth*(`APPRam_depth*0+116)-1:`VWidth*(`APPRam_depth*0+115)]};
			end
			116:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+117)-1:`VWidth*(`APPRam_depth*31+116)],data_in[`VWidth*(`APPRam_depth*30+117)-1:`VWidth*(`APPRam_depth*30+116)],data_in[`VWidth*(`APPRam_depth*29+117)-1:`VWidth*(`APPRam_depth*29+116)],data_in[`VWidth*(`APPRam_depth*28+117)-1:`VWidth*(`APPRam_depth*28+116)],data_in[`VWidth*(`APPRam_depth*27+117)-1:`VWidth*(`APPRam_depth*27+116)],data_in[`VWidth*(`APPRam_depth*26+117)-1:`VWidth*(`APPRam_depth*26+116)],data_in[`VWidth*(`APPRam_depth*25+117)-1:`VWidth*(`APPRam_depth*25+116)],data_in[`VWidth*(`APPRam_depth*24+117)-1:`VWidth*(`APPRam_depth*24+116)],data_in[`VWidth*(`APPRam_depth*23+117)-1:`VWidth*(`APPRam_depth*23+116)],data_in[`VWidth*(`APPRam_depth*22+117)-1:`VWidth*(`APPRam_depth*22+116)],data_in[`VWidth*(`APPRam_depth*21+117)-1:`VWidth*(`APPRam_depth*21+116)],data_in[`VWidth*(`APPRam_depth*20+117)-1:`VWidth*(`APPRam_depth*20+116)],data_in[`VWidth*(`APPRam_depth*19+117)-1:`VWidth*(`APPRam_depth*19+116)],data_in[`VWidth*(`APPRam_depth*18+117)-1:`VWidth*(`APPRam_depth*18+116)],data_in[`VWidth*(`APPRam_depth*17+117)-1:`VWidth*(`APPRam_depth*17+116)],data_in[`VWidth*(`APPRam_depth*16+117)-1:`VWidth*(`APPRam_depth*16+116)],data_in[`VWidth*(`APPRam_depth*15+117)-1:`VWidth*(`APPRam_depth*15+116)],data_in[`VWidth*(`APPRam_depth*14+117)-1:`VWidth*(`APPRam_depth*14+116)],data_in[`VWidth*(`APPRam_depth*13+117)-1:`VWidth*(`APPRam_depth*13+116)],data_in[`VWidth*(`APPRam_depth*12+117)-1:`VWidth*(`APPRam_depth*12+116)],data_in[`VWidth*(`APPRam_depth*11+117)-1:`VWidth*(`APPRam_depth*11+116)],data_in[`VWidth*(`APPRam_depth*10+117)-1:`VWidth*(`APPRam_depth*10+116)],data_in[`VWidth*(`APPRam_depth*9+117)-1:`VWidth*(`APPRam_depth*9+116)],data_in[`VWidth*(`APPRam_depth*8+117)-1:`VWidth*(`APPRam_depth*8+116)],data_in[`VWidth*(`APPRam_depth*7+117)-1:`VWidth*(`APPRam_depth*7+116)],data_in[`VWidth*(`APPRam_depth*6+117)-1:`VWidth*(`APPRam_depth*6+116)],data_in[`VWidth*(`APPRam_depth*5+117)-1:`VWidth*(`APPRam_depth*5+116)],data_in[`VWidth*(`APPRam_depth*4+117)-1:`VWidth*(`APPRam_depth*4+116)],data_in[`VWidth*(`APPRam_depth*3+117)-1:`VWidth*(`APPRam_depth*3+116)],data_in[`VWidth*(`APPRam_depth*2+117)-1:`VWidth*(`APPRam_depth*2+116)],data_in[`VWidth*(`APPRam_depth*1+117)-1:`VWidth*(`APPRam_depth*1+116)],data_in[`VWidth*(`APPRam_depth*0+117)-1:`VWidth*(`APPRam_depth*0+116)]};
			end
			117:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+118)-1:`VWidth*(`APPRam_depth*31+117)],data_in[`VWidth*(`APPRam_depth*30+118)-1:`VWidth*(`APPRam_depth*30+117)],data_in[`VWidth*(`APPRam_depth*29+118)-1:`VWidth*(`APPRam_depth*29+117)],data_in[`VWidth*(`APPRam_depth*28+118)-1:`VWidth*(`APPRam_depth*28+117)],data_in[`VWidth*(`APPRam_depth*27+118)-1:`VWidth*(`APPRam_depth*27+117)],data_in[`VWidth*(`APPRam_depth*26+118)-1:`VWidth*(`APPRam_depth*26+117)],data_in[`VWidth*(`APPRam_depth*25+118)-1:`VWidth*(`APPRam_depth*25+117)],data_in[`VWidth*(`APPRam_depth*24+118)-1:`VWidth*(`APPRam_depth*24+117)],data_in[`VWidth*(`APPRam_depth*23+118)-1:`VWidth*(`APPRam_depth*23+117)],data_in[`VWidth*(`APPRam_depth*22+118)-1:`VWidth*(`APPRam_depth*22+117)],data_in[`VWidth*(`APPRam_depth*21+118)-1:`VWidth*(`APPRam_depth*21+117)],data_in[`VWidth*(`APPRam_depth*20+118)-1:`VWidth*(`APPRam_depth*20+117)],data_in[`VWidth*(`APPRam_depth*19+118)-1:`VWidth*(`APPRam_depth*19+117)],data_in[`VWidth*(`APPRam_depth*18+118)-1:`VWidth*(`APPRam_depth*18+117)],data_in[`VWidth*(`APPRam_depth*17+118)-1:`VWidth*(`APPRam_depth*17+117)],data_in[`VWidth*(`APPRam_depth*16+118)-1:`VWidth*(`APPRam_depth*16+117)],data_in[`VWidth*(`APPRam_depth*15+118)-1:`VWidth*(`APPRam_depth*15+117)],data_in[`VWidth*(`APPRam_depth*14+118)-1:`VWidth*(`APPRam_depth*14+117)],data_in[`VWidth*(`APPRam_depth*13+118)-1:`VWidth*(`APPRam_depth*13+117)],data_in[`VWidth*(`APPRam_depth*12+118)-1:`VWidth*(`APPRam_depth*12+117)],data_in[`VWidth*(`APPRam_depth*11+118)-1:`VWidth*(`APPRam_depth*11+117)],data_in[`VWidth*(`APPRam_depth*10+118)-1:`VWidth*(`APPRam_depth*10+117)],data_in[`VWidth*(`APPRam_depth*9+118)-1:`VWidth*(`APPRam_depth*9+117)],data_in[`VWidth*(`APPRam_depth*8+118)-1:`VWidth*(`APPRam_depth*8+117)],data_in[`VWidth*(`APPRam_depth*7+118)-1:`VWidth*(`APPRam_depth*7+117)],data_in[`VWidth*(`APPRam_depth*6+118)-1:`VWidth*(`APPRam_depth*6+117)],data_in[`VWidth*(`APPRam_depth*5+118)-1:`VWidth*(`APPRam_depth*5+117)],data_in[`VWidth*(`APPRam_depth*4+118)-1:`VWidth*(`APPRam_depth*4+117)],data_in[`VWidth*(`APPRam_depth*3+118)-1:`VWidth*(`APPRam_depth*3+117)],data_in[`VWidth*(`APPRam_depth*2+118)-1:`VWidth*(`APPRam_depth*2+117)],data_in[`VWidth*(`APPRam_depth*1+118)-1:`VWidth*(`APPRam_depth*1+117)],data_in[`VWidth*(`APPRam_depth*0+118)-1:`VWidth*(`APPRam_depth*0+117)]};
			end
			118:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+119)-1:`VWidth*(`APPRam_depth*31+118)],data_in[`VWidth*(`APPRam_depth*30+119)-1:`VWidth*(`APPRam_depth*30+118)],data_in[`VWidth*(`APPRam_depth*29+119)-1:`VWidth*(`APPRam_depth*29+118)],data_in[`VWidth*(`APPRam_depth*28+119)-1:`VWidth*(`APPRam_depth*28+118)],data_in[`VWidth*(`APPRam_depth*27+119)-1:`VWidth*(`APPRam_depth*27+118)],data_in[`VWidth*(`APPRam_depth*26+119)-1:`VWidth*(`APPRam_depth*26+118)],data_in[`VWidth*(`APPRam_depth*25+119)-1:`VWidth*(`APPRam_depth*25+118)],data_in[`VWidth*(`APPRam_depth*24+119)-1:`VWidth*(`APPRam_depth*24+118)],data_in[`VWidth*(`APPRam_depth*23+119)-1:`VWidth*(`APPRam_depth*23+118)],data_in[`VWidth*(`APPRam_depth*22+119)-1:`VWidth*(`APPRam_depth*22+118)],data_in[`VWidth*(`APPRam_depth*21+119)-1:`VWidth*(`APPRam_depth*21+118)],data_in[`VWidth*(`APPRam_depth*20+119)-1:`VWidth*(`APPRam_depth*20+118)],data_in[`VWidth*(`APPRam_depth*19+119)-1:`VWidth*(`APPRam_depth*19+118)],data_in[`VWidth*(`APPRam_depth*18+119)-1:`VWidth*(`APPRam_depth*18+118)],data_in[`VWidth*(`APPRam_depth*17+119)-1:`VWidth*(`APPRam_depth*17+118)],data_in[`VWidth*(`APPRam_depth*16+119)-1:`VWidth*(`APPRam_depth*16+118)],data_in[`VWidth*(`APPRam_depth*15+119)-1:`VWidth*(`APPRam_depth*15+118)],data_in[`VWidth*(`APPRam_depth*14+119)-1:`VWidth*(`APPRam_depth*14+118)],data_in[`VWidth*(`APPRam_depth*13+119)-1:`VWidth*(`APPRam_depth*13+118)],data_in[`VWidth*(`APPRam_depth*12+119)-1:`VWidth*(`APPRam_depth*12+118)],data_in[`VWidth*(`APPRam_depth*11+119)-1:`VWidth*(`APPRam_depth*11+118)],data_in[`VWidth*(`APPRam_depth*10+119)-1:`VWidth*(`APPRam_depth*10+118)],data_in[`VWidth*(`APPRam_depth*9+119)-1:`VWidth*(`APPRam_depth*9+118)],data_in[`VWidth*(`APPRam_depth*8+119)-1:`VWidth*(`APPRam_depth*8+118)],data_in[`VWidth*(`APPRam_depth*7+119)-1:`VWidth*(`APPRam_depth*7+118)],data_in[`VWidth*(`APPRam_depth*6+119)-1:`VWidth*(`APPRam_depth*6+118)],data_in[`VWidth*(`APPRam_depth*5+119)-1:`VWidth*(`APPRam_depth*5+118)],data_in[`VWidth*(`APPRam_depth*4+119)-1:`VWidth*(`APPRam_depth*4+118)],data_in[`VWidth*(`APPRam_depth*3+119)-1:`VWidth*(`APPRam_depth*3+118)],data_in[`VWidth*(`APPRam_depth*2+119)-1:`VWidth*(`APPRam_depth*2+118)],data_in[`VWidth*(`APPRam_depth*1+119)-1:`VWidth*(`APPRam_depth*1+118)],data_in[`VWidth*(`APPRam_depth*0+119)-1:`VWidth*(`APPRam_depth*0+118)]};
			end
			119:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+120)-1:`VWidth*(`APPRam_depth*31+119)],data_in[`VWidth*(`APPRam_depth*30+120)-1:`VWidth*(`APPRam_depth*30+119)],data_in[`VWidth*(`APPRam_depth*29+120)-1:`VWidth*(`APPRam_depth*29+119)],data_in[`VWidth*(`APPRam_depth*28+120)-1:`VWidth*(`APPRam_depth*28+119)],data_in[`VWidth*(`APPRam_depth*27+120)-1:`VWidth*(`APPRam_depth*27+119)],data_in[`VWidth*(`APPRam_depth*26+120)-1:`VWidth*(`APPRam_depth*26+119)],data_in[`VWidth*(`APPRam_depth*25+120)-1:`VWidth*(`APPRam_depth*25+119)],data_in[`VWidth*(`APPRam_depth*24+120)-1:`VWidth*(`APPRam_depth*24+119)],data_in[`VWidth*(`APPRam_depth*23+120)-1:`VWidth*(`APPRam_depth*23+119)],data_in[`VWidth*(`APPRam_depth*22+120)-1:`VWidth*(`APPRam_depth*22+119)],data_in[`VWidth*(`APPRam_depth*21+120)-1:`VWidth*(`APPRam_depth*21+119)],data_in[`VWidth*(`APPRam_depth*20+120)-1:`VWidth*(`APPRam_depth*20+119)],data_in[`VWidth*(`APPRam_depth*19+120)-1:`VWidth*(`APPRam_depth*19+119)],data_in[`VWidth*(`APPRam_depth*18+120)-1:`VWidth*(`APPRam_depth*18+119)],data_in[`VWidth*(`APPRam_depth*17+120)-1:`VWidth*(`APPRam_depth*17+119)],data_in[`VWidth*(`APPRam_depth*16+120)-1:`VWidth*(`APPRam_depth*16+119)],data_in[`VWidth*(`APPRam_depth*15+120)-1:`VWidth*(`APPRam_depth*15+119)],data_in[`VWidth*(`APPRam_depth*14+120)-1:`VWidth*(`APPRam_depth*14+119)],data_in[`VWidth*(`APPRam_depth*13+120)-1:`VWidth*(`APPRam_depth*13+119)],data_in[`VWidth*(`APPRam_depth*12+120)-1:`VWidth*(`APPRam_depth*12+119)],data_in[`VWidth*(`APPRam_depth*11+120)-1:`VWidth*(`APPRam_depth*11+119)],data_in[`VWidth*(`APPRam_depth*10+120)-1:`VWidth*(`APPRam_depth*10+119)],data_in[`VWidth*(`APPRam_depth*9+120)-1:`VWidth*(`APPRam_depth*9+119)],data_in[`VWidth*(`APPRam_depth*8+120)-1:`VWidth*(`APPRam_depth*8+119)],data_in[`VWidth*(`APPRam_depth*7+120)-1:`VWidth*(`APPRam_depth*7+119)],data_in[`VWidth*(`APPRam_depth*6+120)-1:`VWidth*(`APPRam_depth*6+119)],data_in[`VWidth*(`APPRam_depth*5+120)-1:`VWidth*(`APPRam_depth*5+119)],data_in[`VWidth*(`APPRam_depth*4+120)-1:`VWidth*(`APPRam_depth*4+119)],data_in[`VWidth*(`APPRam_depth*3+120)-1:`VWidth*(`APPRam_depth*3+119)],data_in[`VWidth*(`APPRam_depth*2+120)-1:`VWidth*(`APPRam_depth*2+119)],data_in[`VWidth*(`APPRam_depth*1+120)-1:`VWidth*(`APPRam_depth*1+119)],data_in[`VWidth*(`APPRam_depth*0+120)-1:`VWidth*(`APPRam_depth*0+119)]};
			end
			120:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+121)-1:`VWidth*(`APPRam_depth*31+120)],data_in[`VWidth*(`APPRam_depth*30+121)-1:`VWidth*(`APPRam_depth*30+120)],data_in[`VWidth*(`APPRam_depth*29+121)-1:`VWidth*(`APPRam_depth*29+120)],data_in[`VWidth*(`APPRam_depth*28+121)-1:`VWidth*(`APPRam_depth*28+120)],data_in[`VWidth*(`APPRam_depth*27+121)-1:`VWidth*(`APPRam_depth*27+120)],data_in[`VWidth*(`APPRam_depth*26+121)-1:`VWidth*(`APPRam_depth*26+120)],data_in[`VWidth*(`APPRam_depth*25+121)-1:`VWidth*(`APPRam_depth*25+120)],data_in[`VWidth*(`APPRam_depth*24+121)-1:`VWidth*(`APPRam_depth*24+120)],data_in[`VWidth*(`APPRam_depth*23+121)-1:`VWidth*(`APPRam_depth*23+120)],data_in[`VWidth*(`APPRam_depth*22+121)-1:`VWidth*(`APPRam_depth*22+120)],data_in[`VWidth*(`APPRam_depth*21+121)-1:`VWidth*(`APPRam_depth*21+120)],data_in[`VWidth*(`APPRam_depth*20+121)-1:`VWidth*(`APPRam_depth*20+120)],data_in[`VWidth*(`APPRam_depth*19+121)-1:`VWidth*(`APPRam_depth*19+120)],data_in[`VWidth*(`APPRam_depth*18+121)-1:`VWidth*(`APPRam_depth*18+120)],data_in[`VWidth*(`APPRam_depth*17+121)-1:`VWidth*(`APPRam_depth*17+120)],data_in[`VWidth*(`APPRam_depth*16+121)-1:`VWidth*(`APPRam_depth*16+120)],data_in[`VWidth*(`APPRam_depth*15+121)-1:`VWidth*(`APPRam_depth*15+120)],data_in[`VWidth*(`APPRam_depth*14+121)-1:`VWidth*(`APPRam_depth*14+120)],data_in[`VWidth*(`APPRam_depth*13+121)-1:`VWidth*(`APPRam_depth*13+120)],data_in[`VWidth*(`APPRam_depth*12+121)-1:`VWidth*(`APPRam_depth*12+120)],data_in[`VWidth*(`APPRam_depth*11+121)-1:`VWidth*(`APPRam_depth*11+120)],data_in[`VWidth*(`APPRam_depth*10+121)-1:`VWidth*(`APPRam_depth*10+120)],data_in[`VWidth*(`APPRam_depth*9+121)-1:`VWidth*(`APPRam_depth*9+120)],data_in[`VWidth*(`APPRam_depth*8+121)-1:`VWidth*(`APPRam_depth*8+120)],data_in[`VWidth*(`APPRam_depth*7+121)-1:`VWidth*(`APPRam_depth*7+120)],data_in[`VWidth*(`APPRam_depth*6+121)-1:`VWidth*(`APPRam_depth*6+120)],data_in[`VWidth*(`APPRam_depth*5+121)-1:`VWidth*(`APPRam_depth*5+120)],data_in[`VWidth*(`APPRam_depth*4+121)-1:`VWidth*(`APPRam_depth*4+120)],data_in[`VWidth*(`APPRam_depth*3+121)-1:`VWidth*(`APPRam_depth*3+120)],data_in[`VWidth*(`APPRam_depth*2+121)-1:`VWidth*(`APPRam_depth*2+120)],data_in[`VWidth*(`APPRam_depth*1+121)-1:`VWidth*(`APPRam_depth*1+120)],data_in[`VWidth*(`APPRam_depth*0+121)-1:`VWidth*(`APPRam_depth*0+120)]};
			end
			121:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+122)-1:`VWidth*(`APPRam_depth*31+121)],data_in[`VWidth*(`APPRam_depth*30+122)-1:`VWidth*(`APPRam_depth*30+121)],data_in[`VWidth*(`APPRam_depth*29+122)-1:`VWidth*(`APPRam_depth*29+121)],data_in[`VWidth*(`APPRam_depth*28+122)-1:`VWidth*(`APPRam_depth*28+121)],data_in[`VWidth*(`APPRam_depth*27+122)-1:`VWidth*(`APPRam_depth*27+121)],data_in[`VWidth*(`APPRam_depth*26+122)-1:`VWidth*(`APPRam_depth*26+121)],data_in[`VWidth*(`APPRam_depth*25+122)-1:`VWidth*(`APPRam_depth*25+121)],data_in[`VWidth*(`APPRam_depth*24+122)-1:`VWidth*(`APPRam_depth*24+121)],data_in[`VWidth*(`APPRam_depth*23+122)-1:`VWidth*(`APPRam_depth*23+121)],data_in[`VWidth*(`APPRam_depth*22+122)-1:`VWidth*(`APPRam_depth*22+121)],data_in[`VWidth*(`APPRam_depth*21+122)-1:`VWidth*(`APPRam_depth*21+121)],data_in[`VWidth*(`APPRam_depth*20+122)-1:`VWidth*(`APPRam_depth*20+121)],data_in[`VWidth*(`APPRam_depth*19+122)-1:`VWidth*(`APPRam_depth*19+121)],data_in[`VWidth*(`APPRam_depth*18+122)-1:`VWidth*(`APPRam_depth*18+121)],data_in[`VWidth*(`APPRam_depth*17+122)-1:`VWidth*(`APPRam_depth*17+121)],data_in[`VWidth*(`APPRam_depth*16+122)-1:`VWidth*(`APPRam_depth*16+121)],data_in[`VWidth*(`APPRam_depth*15+122)-1:`VWidth*(`APPRam_depth*15+121)],data_in[`VWidth*(`APPRam_depth*14+122)-1:`VWidth*(`APPRam_depth*14+121)],data_in[`VWidth*(`APPRam_depth*13+122)-1:`VWidth*(`APPRam_depth*13+121)],data_in[`VWidth*(`APPRam_depth*12+122)-1:`VWidth*(`APPRam_depth*12+121)],data_in[`VWidth*(`APPRam_depth*11+122)-1:`VWidth*(`APPRam_depth*11+121)],data_in[`VWidth*(`APPRam_depth*10+122)-1:`VWidth*(`APPRam_depth*10+121)],data_in[`VWidth*(`APPRam_depth*9+122)-1:`VWidth*(`APPRam_depth*9+121)],data_in[`VWidth*(`APPRam_depth*8+122)-1:`VWidth*(`APPRam_depth*8+121)],data_in[`VWidth*(`APPRam_depth*7+122)-1:`VWidth*(`APPRam_depth*7+121)],data_in[`VWidth*(`APPRam_depth*6+122)-1:`VWidth*(`APPRam_depth*6+121)],data_in[`VWidth*(`APPRam_depth*5+122)-1:`VWidth*(`APPRam_depth*5+121)],data_in[`VWidth*(`APPRam_depth*4+122)-1:`VWidth*(`APPRam_depth*4+121)],data_in[`VWidth*(`APPRam_depth*3+122)-1:`VWidth*(`APPRam_depth*3+121)],data_in[`VWidth*(`APPRam_depth*2+122)-1:`VWidth*(`APPRam_depth*2+121)],data_in[`VWidth*(`APPRam_depth*1+122)-1:`VWidth*(`APPRam_depth*1+121)],data_in[`VWidth*(`APPRam_depth*0+122)-1:`VWidth*(`APPRam_depth*0+121)]};
			end
			122:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+123)-1:`VWidth*(`APPRam_depth*31+122)],data_in[`VWidth*(`APPRam_depth*30+123)-1:`VWidth*(`APPRam_depth*30+122)],data_in[`VWidth*(`APPRam_depth*29+123)-1:`VWidth*(`APPRam_depth*29+122)],data_in[`VWidth*(`APPRam_depth*28+123)-1:`VWidth*(`APPRam_depth*28+122)],data_in[`VWidth*(`APPRam_depth*27+123)-1:`VWidth*(`APPRam_depth*27+122)],data_in[`VWidth*(`APPRam_depth*26+123)-1:`VWidth*(`APPRam_depth*26+122)],data_in[`VWidth*(`APPRam_depth*25+123)-1:`VWidth*(`APPRam_depth*25+122)],data_in[`VWidth*(`APPRam_depth*24+123)-1:`VWidth*(`APPRam_depth*24+122)],data_in[`VWidth*(`APPRam_depth*23+123)-1:`VWidth*(`APPRam_depth*23+122)],data_in[`VWidth*(`APPRam_depth*22+123)-1:`VWidth*(`APPRam_depth*22+122)],data_in[`VWidth*(`APPRam_depth*21+123)-1:`VWidth*(`APPRam_depth*21+122)],data_in[`VWidth*(`APPRam_depth*20+123)-1:`VWidth*(`APPRam_depth*20+122)],data_in[`VWidth*(`APPRam_depth*19+123)-1:`VWidth*(`APPRam_depth*19+122)],data_in[`VWidth*(`APPRam_depth*18+123)-1:`VWidth*(`APPRam_depth*18+122)],data_in[`VWidth*(`APPRam_depth*17+123)-1:`VWidth*(`APPRam_depth*17+122)],data_in[`VWidth*(`APPRam_depth*16+123)-1:`VWidth*(`APPRam_depth*16+122)],data_in[`VWidth*(`APPRam_depth*15+123)-1:`VWidth*(`APPRam_depth*15+122)],data_in[`VWidth*(`APPRam_depth*14+123)-1:`VWidth*(`APPRam_depth*14+122)],data_in[`VWidth*(`APPRam_depth*13+123)-1:`VWidth*(`APPRam_depth*13+122)],data_in[`VWidth*(`APPRam_depth*12+123)-1:`VWidth*(`APPRam_depth*12+122)],data_in[`VWidth*(`APPRam_depth*11+123)-1:`VWidth*(`APPRam_depth*11+122)],data_in[`VWidth*(`APPRam_depth*10+123)-1:`VWidth*(`APPRam_depth*10+122)],data_in[`VWidth*(`APPRam_depth*9+123)-1:`VWidth*(`APPRam_depth*9+122)],data_in[`VWidth*(`APPRam_depth*8+123)-1:`VWidth*(`APPRam_depth*8+122)],data_in[`VWidth*(`APPRam_depth*7+123)-1:`VWidth*(`APPRam_depth*7+122)],data_in[`VWidth*(`APPRam_depth*6+123)-1:`VWidth*(`APPRam_depth*6+122)],data_in[`VWidth*(`APPRam_depth*5+123)-1:`VWidth*(`APPRam_depth*5+122)],data_in[`VWidth*(`APPRam_depth*4+123)-1:`VWidth*(`APPRam_depth*4+122)],data_in[`VWidth*(`APPRam_depth*3+123)-1:`VWidth*(`APPRam_depth*3+122)],data_in[`VWidth*(`APPRam_depth*2+123)-1:`VWidth*(`APPRam_depth*2+122)],data_in[`VWidth*(`APPRam_depth*1+123)-1:`VWidth*(`APPRam_depth*1+122)],data_in[`VWidth*(`APPRam_depth*0+123)-1:`VWidth*(`APPRam_depth*0+122)]};
			end
			123:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+124)-1:`VWidth*(`APPRam_depth*31+123)],data_in[`VWidth*(`APPRam_depth*30+124)-1:`VWidth*(`APPRam_depth*30+123)],data_in[`VWidth*(`APPRam_depth*29+124)-1:`VWidth*(`APPRam_depth*29+123)],data_in[`VWidth*(`APPRam_depth*28+124)-1:`VWidth*(`APPRam_depth*28+123)],data_in[`VWidth*(`APPRam_depth*27+124)-1:`VWidth*(`APPRam_depth*27+123)],data_in[`VWidth*(`APPRam_depth*26+124)-1:`VWidth*(`APPRam_depth*26+123)],data_in[`VWidth*(`APPRam_depth*25+124)-1:`VWidth*(`APPRam_depth*25+123)],data_in[`VWidth*(`APPRam_depth*24+124)-1:`VWidth*(`APPRam_depth*24+123)],data_in[`VWidth*(`APPRam_depth*23+124)-1:`VWidth*(`APPRam_depth*23+123)],data_in[`VWidth*(`APPRam_depth*22+124)-1:`VWidth*(`APPRam_depth*22+123)],data_in[`VWidth*(`APPRam_depth*21+124)-1:`VWidth*(`APPRam_depth*21+123)],data_in[`VWidth*(`APPRam_depth*20+124)-1:`VWidth*(`APPRam_depth*20+123)],data_in[`VWidth*(`APPRam_depth*19+124)-1:`VWidth*(`APPRam_depth*19+123)],data_in[`VWidth*(`APPRam_depth*18+124)-1:`VWidth*(`APPRam_depth*18+123)],data_in[`VWidth*(`APPRam_depth*17+124)-1:`VWidth*(`APPRam_depth*17+123)],data_in[`VWidth*(`APPRam_depth*16+124)-1:`VWidth*(`APPRam_depth*16+123)],data_in[`VWidth*(`APPRam_depth*15+124)-1:`VWidth*(`APPRam_depth*15+123)],data_in[`VWidth*(`APPRam_depth*14+124)-1:`VWidth*(`APPRam_depth*14+123)],data_in[`VWidth*(`APPRam_depth*13+124)-1:`VWidth*(`APPRam_depth*13+123)],data_in[`VWidth*(`APPRam_depth*12+124)-1:`VWidth*(`APPRam_depth*12+123)],data_in[`VWidth*(`APPRam_depth*11+124)-1:`VWidth*(`APPRam_depth*11+123)],data_in[`VWidth*(`APPRam_depth*10+124)-1:`VWidth*(`APPRam_depth*10+123)],data_in[`VWidth*(`APPRam_depth*9+124)-1:`VWidth*(`APPRam_depth*9+123)],data_in[`VWidth*(`APPRam_depth*8+124)-1:`VWidth*(`APPRam_depth*8+123)],data_in[`VWidth*(`APPRam_depth*7+124)-1:`VWidth*(`APPRam_depth*7+123)],data_in[`VWidth*(`APPRam_depth*6+124)-1:`VWidth*(`APPRam_depth*6+123)],data_in[`VWidth*(`APPRam_depth*5+124)-1:`VWidth*(`APPRam_depth*5+123)],data_in[`VWidth*(`APPRam_depth*4+124)-1:`VWidth*(`APPRam_depth*4+123)],data_in[`VWidth*(`APPRam_depth*3+124)-1:`VWidth*(`APPRam_depth*3+123)],data_in[`VWidth*(`APPRam_depth*2+124)-1:`VWidth*(`APPRam_depth*2+123)],data_in[`VWidth*(`APPRam_depth*1+124)-1:`VWidth*(`APPRam_depth*1+123)],data_in[`VWidth*(`APPRam_depth*0+124)-1:`VWidth*(`APPRam_depth*0+123)]};
			end
			124:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+125)-1:`VWidth*(`APPRam_depth*31+124)],data_in[`VWidth*(`APPRam_depth*30+125)-1:`VWidth*(`APPRam_depth*30+124)],data_in[`VWidth*(`APPRam_depth*29+125)-1:`VWidth*(`APPRam_depth*29+124)],data_in[`VWidth*(`APPRam_depth*28+125)-1:`VWidth*(`APPRam_depth*28+124)],data_in[`VWidth*(`APPRam_depth*27+125)-1:`VWidth*(`APPRam_depth*27+124)],data_in[`VWidth*(`APPRam_depth*26+125)-1:`VWidth*(`APPRam_depth*26+124)],data_in[`VWidth*(`APPRam_depth*25+125)-1:`VWidth*(`APPRam_depth*25+124)],data_in[`VWidth*(`APPRam_depth*24+125)-1:`VWidth*(`APPRam_depth*24+124)],data_in[`VWidth*(`APPRam_depth*23+125)-1:`VWidth*(`APPRam_depth*23+124)],data_in[`VWidth*(`APPRam_depth*22+125)-1:`VWidth*(`APPRam_depth*22+124)],data_in[`VWidth*(`APPRam_depth*21+125)-1:`VWidth*(`APPRam_depth*21+124)],data_in[`VWidth*(`APPRam_depth*20+125)-1:`VWidth*(`APPRam_depth*20+124)],data_in[`VWidth*(`APPRam_depth*19+125)-1:`VWidth*(`APPRam_depth*19+124)],data_in[`VWidth*(`APPRam_depth*18+125)-1:`VWidth*(`APPRam_depth*18+124)],data_in[`VWidth*(`APPRam_depth*17+125)-1:`VWidth*(`APPRam_depth*17+124)],data_in[`VWidth*(`APPRam_depth*16+125)-1:`VWidth*(`APPRam_depth*16+124)],data_in[`VWidth*(`APPRam_depth*15+125)-1:`VWidth*(`APPRam_depth*15+124)],data_in[`VWidth*(`APPRam_depth*14+125)-1:`VWidth*(`APPRam_depth*14+124)],data_in[`VWidth*(`APPRam_depth*13+125)-1:`VWidth*(`APPRam_depth*13+124)],data_in[`VWidth*(`APPRam_depth*12+125)-1:`VWidth*(`APPRam_depth*12+124)],data_in[`VWidth*(`APPRam_depth*11+125)-1:`VWidth*(`APPRam_depth*11+124)],data_in[`VWidth*(`APPRam_depth*10+125)-1:`VWidth*(`APPRam_depth*10+124)],data_in[`VWidth*(`APPRam_depth*9+125)-1:`VWidth*(`APPRam_depth*9+124)],data_in[`VWidth*(`APPRam_depth*8+125)-1:`VWidth*(`APPRam_depth*8+124)],data_in[`VWidth*(`APPRam_depth*7+125)-1:`VWidth*(`APPRam_depth*7+124)],data_in[`VWidth*(`APPRam_depth*6+125)-1:`VWidth*(`APPRam_depth*6+124)],data_in[`VWidth*(`APPRam_depth*5+125)-1:`VWidth*(`APPRam_depth*5+124)],data_in[`VWidth*(`APPRam_depth*4+125)-1:`VWidth*(`APPRam_depth*4+124)],data_in[`VWidth*(`APPRam_depth*3+125)-1:`VWidth*(`APPRam_depth*3+124)],data_in[`VWidth*(`APPRam_depth*2+125)-1:`VWidth*(`APPRam_depth*2+124)],data_in[`VWidth*(`APPRam_depth*1+125)-1:`VWidth*(`APPRam_depth*1+124)],data_in[`VWidth*(`APPRam_depth*0+125)-1:`VWidth*(`APPRam_depth*0+124)]};
			end
			125:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+126)-1:`VWidth*(`APPRam_depth*31+125)],data_in[`VWidth*(`APPRam_depth*30+126)-1:`VWidth*(`APPRam_depth*30+125)],data_in[`VWidth*(`APPRam_depth*29+126)-1:`VWidth*(`APPRam_depth*29+125)],data_in[`VWidth*(`APPRam_depth*28+126)-1:`VWidth*(`APPRam_depth*28+125)],data_in[`VWidth*(`APPRam_depth*27+126)-1:`VWidth*(`APPRam_depth*27+125)],data_in[`VWidth*(`APPRam_depth*26+126)-1:`VWidth*(`APPRam_depth*26+125)],data_in[`VWidth*(`APPRam_depth*25+126)-1:`VWidth*(`APPRam_depth*25+125)],data_in[`VWidth*(`APPRam_depth*24+126)-1:`VWidth*(`APPRam_depth*24+125)],data_in[`VWidth*(`APPRam_depth*23+126)-1:`VWidth*(`APPRam_depth*23+125)],data_in[`VWidth*(`APPRam_depth*22+126)-1:`VWidth*(`APPRam_depth*22+125)],data_in[`VWidth*(`APPRam_depth*21+126)-1:`VWidth*(`APPRam_depth*21+125)],data_in[`VWidth*(`APPRam_depth*20+126)-1:`VWidth*(`APPRam_depth*20+125)],data_in[`VWidth*(`APPRam_depth*19+126)-1:`VWidth*(`APPRam_depth*19+125)],data_in[`VWidth*(`APPRam_depth*18+126)-1:`VWidth*(`APPRam_depth*18+125)],data_in[`VWidth*(`APPRam_depth*17+126)-1:`VWidth*(`APPRam_depth*17+125)],data_in[`VWidth*(`APPRam_depth*16+126)-1:`VWidth*(`APPRam_depth*16+125)],data_in[`VWidth*(`APPRam_depth*15+126)-1:`VWidth*(`APPRam_depth*15+125)],data_in[`VWidth*(`APPRam_depth*14+126)-1:`VWidth*(`APPRam_depth*14+125)],data_in[`VWidth*(`APPRam_depth*13+126)-1:`VWidth*(`APPRam_depth*13+125)],data_in[`VWidth*(`APPRam_depth*12+126)-1:`VWidth*(`APPRam_depth*12+125)],data_in[`VWidth*(`APPRam_depth*11+126)-1:`VWidth*(`APPRam_depth*11+125)],data_in[`VWidth*(`APPRam_depth*10+126)-1:`VWidth*(`APPRam_depth*10+125)],data_in[`VWidth*(`APPRam_depth*9+126)-1:`VWidth*(`APPRam_depth*9+125)],data_in[`VWidth*(`APPRam_depth*8+126)-1:`VWidth*(`APPRam_depth*8+125)],data_in[`VWidth*(`APPRam_depth*7+126)-1:`VWidth*(`APPRam_depth*7+125)],data_in[`VWidth*(`APPRam_depth*6+126)-1:`VWidth*(`APPRam_depth*6+125)],data_in[`VWidth*(`APPRam_depth*5+126)-1:`VWidth*(`APPRam_depth*5+125)],data_in[`VWidth*(`APPRam_depth*4+126)-1:`VWidth*(`APPRam_depth*4+125)],data_in[`VWidth*(`APPRam_depth*3+126)-1:`VWidth*(`APPRam_depth*3+125)],data_in[`VWidth*(`APPRam_depth*2+126)-1:`VWidth*(`APPRam_depth*2+125)],data_in[`VWidth*(`APPRam_depth*1+126)-1:`VWidth*(`APPRam_depth*1+125)],data_in[`VWidth*(`APPRam_depth*0+126)-1:`VWidth*(`APPRam_depth*0+125)]};
			end
			126:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+127)-1:`VWidth*(`APPRam_depth*31+126)],data_in[`VWidth*(`APPRam_depth*30+127)-1:`VWidth*(`APPRam_depth*30+126)],data_in[`VWidth*(`APPRam_depth*29+127)-1:`VWidth*(`APPRam_depth*29+126)],data_in[`VWidth*(`APPRam_depth*28+127)-1:`VWidth*(`APPRam_depth*28+126)],data_in[`VWidth*(`APPRam_depth*27+127)-1:`VWidth*(`APPRam_depth*27+126)],data_in[`VWidth*(`APPRam_depth*26+127)-1:`VWidth*(`APPRam_depth*26+126)],data_in[`VWidth*(`APPRam_depth*25+127)-1:`VWidth*(`APPRam_depth*25+126)],data_in[`VWidth*(`APPRam_depth*24+127)-1:`VWidth*(`APPRam_depth*24+126)],data_in[`VWidth*(`APPRam_depth*23+127)-1:`VWidth*(`APPRam_depth*23+126)],data_in[`VWidth*(`APPRam_depth*22+127)-1:`VWidth*(`APPRam_depth*22+126)],data_in[`VWidth*(`APPRam_depth*21+127)-1:`VWidth*(`APPRam_depth*21+126)],data_in[`VWidth*(`APPRam_depth*20+127)-1:`VWidth*(`APPRam_depth*20+126)],data_in[`VWidth*(`APPRam_depth*19+127)-1:`VWidth*(`APPRam_depth*19+126)],data_in[`VWidth*(`APPRam_depth*18+127)-1:`VWidth*(`APPRam_depth*18+126)],data_in[`VWidth*(`APPRam_depth*17+127)-1:`VWidth*(`APPRam_depth*17+126)],data_in[`VWidth*(`APPRam_depth*16+127)-1:`VWidth*(`APPRam_depth*16+126)],data_in[`VWidth*(`APPRam_depth*15+127)-1:`VWidth*(`APPRam_depth*15+126)],data_in[`VWidth*(`APPRam_depth*14+127)-1:`VWidth*(`APPRam_depth*14+126)],data_in[`VWidth*(`APPRam_depth*13+127)-1:`VWidth*(`APPRam_depth*13+126)],data_in[`VWidth*(`APPRam_depth*12+127)-1:`VWidth*(`APPRam_depth*12+126)],data_in[`VWidth*(`APPRam_depth*11+127)-1:`VWidth*(`APPRam_depth*11+126)],data_in[`VWidth*(`APPRam_depth*10+127)-1:`VWidth*(`APPRam_depth*10+126)],data_in[`VWidth*(`APPRam_depth*9+127)-1:`VWidth*(`APPRam_depth*9+126)],data_in[`VWidth*(`APPRam_depth*8+127)-1:`VWidth*(`APPRam_depth*8+126)],data_in[`VWidth*(`APPRam_depth*7+127)-1:`VWidth*(`APPRam_depth*7+126)],data_in[`VWidth*(`APPRam_depth*6+127)-1:`VWidth*(`APPRam_depth*6+126)],data_in[`VWidth*(`APPRam_depth*5+127)-1:`VWidth*(`APPRam_depth*5+126)],data_in[`VWidth*(`APPRam_depth*4+127)-1:`VWidth*(`APPRam_depth*4+126)],data_in[`VWidth*(`APPRam_depth*3+127)-1:`VWidth*(`APPRam_depth*3+126)],data_in[`VWidth*(`APPRam_depth*2+127)-1:`VWidth*(`APPRam_depth*2+126)],data_in[`VWidth*(`APPRam_depth*1+127)-1:`VWidth*(`APPRam_depth*1+126)],data_in[`VWidth*(`APPRam_depth*0+127)-1:`VWidth*(`APPRam_depth*0+126)]};
			end
			127:
			begin
				data_out = {data_in[`VWidth*(`APPRam_depth*31+128)-1:`VWidth*(`APPRam_depth*31+127)],data_in[`VWidth*(`APPRam_depth*30+128)-1:`VWidth*(`APPRam_depth*30+127)],data_in[`VWidth*(`APPRam_depth*29+128)-1:`VWidth*(`APPRam_depth*29+127)],data_in[`VWidth*(`APPRam_depth*28+128)-1:`VWidth*(`APPRam_depth*28+127)],data_in[`VWidth*(`APPRam_depth*27+128)-1:`VWidth*(`APPRam_depth*27+127)],data_in[`VWidth*(`APPRam_depth*26+128)-1:`VWidth*(`APPRam_depth*26+127)],data_in[`VWidth*(`APPRam_depth*25+128)-1:`VWidth*(`APPRam_depth*25+127)],data_in[`VWidth*(`APPRam_depth*24+128)-1:`VWidth*(`APPRam_depth*24+127)],data_in[`VWidth*(`APPRam_depth*23+128)-1:`VWidth*(`APPRam_depth*23+127)],data_in[`VWidth*(`APPRam_depth*22+128)-1:`VWidth*(`APPRam_depth*22+127)],data_in[`VWidth*(`APPRam_depth*21+128)-1:`VWidth*(`APPRam_depth*21+127)],data_in[`VWidth*(`APPRam_depth*20+128)-1:`VWidth*(`APPRam_depth*20+127)],data_in[`VWidth*(`APPRam_depth*19+128)-1:`VWidth*(`APPRam_depth*19+127)],data_in[`VWidth*(`APPRam_depth*18+128)-1:`VWidth*(`APPRam_depth*18+127)],data_in[`VWidth*(`APPRam_depth*17+128)-1:`VWidth*(`APPRam_depth*17+127)],data_in[`VWidth*(`APPRam_depth*16+128)-1:`VWidth*(`APPRam_depth*16+127)],data_in[`VWidth*(`APPRam_depth*15+128)-1:`VWidth*(`APPRam_depth*15+127)],data_in[`VWidth*(`APPRam_depth*14+128)-1:`VWidth*(`APPRam_depth*14+127)],data_in[`VWidth*(`APPRam_depth*13+128)-1:`VWidth*(`APPRam_depth*13+127)],data_in[`VWidth*(`APPRam_depth*12+128)-1:`VWidth*(`APPRam_depth*12+127)],data_in[`VWidth*(`APPRam_depth*11+128)-1:`VWidth*(`APPRam_depth*11+127)],data_in[`VWidth*(`APPRam_depth*10+128)-1:`VWidth*(`APPRam_depth*10+127)],data_in[`VWidth*(`APPRam_depth*9+128)-1:`VWidth*(`APPRam_depth*9+127)],data_in[`VWidth*(`APPRam_depth*8+128)-1:`VWidth*(`APPRam_depth*8+127)],data_in[`VWidth*(`APPRam_depth*7+128)-1:`VWidth*(`APPRam_depth*7+127)],data_in[`VWidth*(`APPRam_depth*6+128)-1:`VWidth*(`APPRam_depth*6+127)],data_in[`VWidth*(`APPRam_depth*5+128)-1:`VWidth*(`APPRam_depth*5+127)],data_in[`VWidth*(`APPRam_depth*4+128)-1:`VWidth*(`APPRam_depth*4+127)],data_in[`VWidth*(`APPRam_depth*3+128)-1:`VWidth*(`APPRam_depth*3+127)],data_in[`VWidth*(`APPRam_depth*2+128)-1:`VWidth*(`APPRam_depth*2+127)],data_in[`VWidth*(`APPRam_depth*1+128)-1:`VWidth*(`APPRam_depth*1+127)],data_in[`VWidth*(`APPRam_depth*0+128)-1:`VWidth*(`APPRam_depth*0+127)]};
			end

			default:
			begin
				data_out <= 0;
			end
		endcase
	end
	else
	begin
		data_out <= 0;
	end
end


endmodule